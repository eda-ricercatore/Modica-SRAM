* Andrew Mattheisen amattheisen@yahoo.com
* Zhiyang Ong zhiyang@ieee.org
* # FILE NAME: /HOME/SCF-08/MATTHEIS/SIMULATION/SRAM_128X256BIT_TOP/HSPICES/    
* SCHEMATIC/NETLIST/SRAM_128X256BIT_TOP.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON OCT 25 01:12:31 2007
   
* GLOBAL NET DEFINITIONS
.GLOBAL VDD! 
* FILE NAME: SRAM2_SRAM_128X256BIT_TOP_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SRAM_128X256BIT_TOP.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:43 2007.
   
XI101 NET0104_0 NET0104_1 NET0104_2 NET0104_3 NET0104_4 NET0104_5 NET0104_6 
+ADDRESS_A_0 ADDRESS_A_1 ADDRESS_A_2 ADDRESS_A_3 ADDRESS_A_4 ADDRESS_A_5 
+ADDRESS_A_6 TL_PI_MODEL7_G13 
XI99 NET0105_0 NET0105_1 NET0105_2 ADDRESS_A_7 ADDRESS_A_8 ADDRESS_A_9 
+TL_PI_MODEL3_G14 
XI95 WRITE_EN_FF WRITE_EN_REAL TL_PI_MODEL_1 
XI98 NET130 CLK TL_PI_MODEL_2 
XI94 NET262_0 NET262_1 NET262_2 NET262_3 NET262_4 NET262_5 NET262_6 NET262_7 
+NET262_8 NET262_9 NET262_10 NET262_11 NET262_12 NET262_13 NET262_14 NET262_15 
+NET262_16 NET262_17 NET262_18 NET262_19 NET262_20 NET262_21 NET262_22 
+NET262_23 NET262_24 NET262_25 NET262_26 NET262_27 NET262_28 NET262_29 
+NET262_30 NET262_31 NET112_0 NET112_1 NET112_2 NET112_3 NET112_4 NET112_5 
+NET112_6 NET112_7 NET112_8 NET112_9 NET112_10 NET112_11 NET112_12 NET112_13 
+NET112_14 NET112_15 NET112_16 NET112_17 NET112_18 NET112_19 NET112_20 
+NET112_21 NET112_22 NET112_23 NET112_24 NET112_25 NET112_26 NET112_27 
+NET112_28 NET112_29 NET112_30 NET112_31 TL_PI_MODEL32_3 
XI92 NET257_0 NET257_1 NET257_2 NET257_3 NET257_4 NET257_5 NET257_6 NET257_7 
+NET257_8 NET257_9 NET257_10 NET257_11 NET257_12 NET257_13 NET257_14 NET257_15 
+NET257_16 NET257_17 NET257_18 NET257_19 NET257_20 NET257_21 NET257_22 
+NET257_23 NET257_24 NET257_25 NET257_26 NET257_27 NET257_28 NET257_29 
+NET257_30 NET257_31 OUT_B_PRE_FF_0 OUT_B_PRE_FF_1 OUT_B_PRE_FF_2 
+OUT_B_PRE_FF_3 OUT_B_PRE_FF_4 OUT_B_PRE_FF_5 OUT_B_PRE_FF_6 OUT_B_PRE_FF_7 
+OUT_B_PRE_FF_8 OUT_B_PRE_FF_9 OUT_B_PRE_FF_10 OUT_B_PRE_FF_11 OUT_B_PRE_FF_12 
+OUT_B_PRE_FF_13 OUT_B_PRE_FF_14 OUT_B_PRE_FF_15 OUT_B_PRE_FF_16 
+OUT_B_PRE_FF_17 OUT_B_PRE_FF_18 OUT_B_PRE_FF_19 OUT_B_PRE_FF_20 
+OUT_B_PRE_FF_21 OUT_B_PRE_FF_22 OUT_B_PRE_FF_23 OUT_B_PRE_FF_24 
+OUT_B_PRE_FF_25 OUT_B_PRE_FF_26 OUT_B_PRE_FF_27 OUT_B_PRE_FF_28 
+OUT_B_PRE_FF_29 OUT_B_PRE_FF_30 OUT_B_PRE_FF_31 TL_PI_MODEL32_4 
XI93 NET260_0 NET260_1 NET260_2 NET260_3 NET260_4 NET260_5 NET260_6 NET260_7 
+NET260_8 NET260_9 NET260_10 NET260_11 NET260_12 NET260_13 NET260_14 NET260_15 
+NET260_16 NET260_17 NET260_18 NET260_19 NET260_20 NET260_21 NET260_22 
+NET260_23 NET260_24 NET260_25 NET260_26 NET260_27 NET260_28 NET260_29 
+NET260_30 NET260_31 NET116_0 NET116_1 NET116_2 NET116_3 NET116_4 NET116_5 
+NET116_6 NET116_7 NET116_8 NET116_9 NET116_10 NET116_11 NET116_12 NET116_13 
+NET116_14 NET116_15 NET116_16 NET116_17 NET116_18 NET116_19 NET116_20 
+NET116_21 NET116_22 NET116_23 NET116_24 NET116_25 NET116_26 NET116_27 
+NET116_28 NET116_29 NET116_30 NET116_31 TL_PI_MODEL32_4 
XI90 CLK WRITE_EN WRITE_EN_FF DFFPOSX1_G6 
XPRECONTROL CLK PRE_REAL READ_EN_REAL WORD_EN_REAL WRITE_EN_REAL DUMMY_ROW_G15 
XI76 NET126 NET124 CLKBUF3_G16 
XI77 NET128 NET126 CLKBUF3_G16 
XI78 CLK_RAW NET128 CLKBUF3_G16 
XI97 NET124 NET130 CLKBUF3_G16 
XI72 NET220_0 NET220_1 NET220_2 NET220_3 NET220_4 NET220_5 NET220_6 NET220_7 
+NET220_8 NET220_9 NET220_10 NET220_11 NET220_12 NET220_13 NET220_14 NET220_15 
+NET220_16 NET220_17 NET220_18 NET220_19 NET220_20 NET220_21 NET220_22 
+NET220_23 NET220_24 NET220_25 NET220_26 NET220_27 NET220_28 NET220_29 
+NET220_30 NET220_31 NET133_0 NET133_1 NET133_2 NET133_3 NET133_4 NET133_5 
+NET133_6 NET133_7 NET133_8 NET133_9 NET133_10 NET133_11 NET133_12 NET133_13 
+NET133_14 NET133_15 NET133_16 NET133_17 NET133_18 NET133_19 NET133_20 
+NET133_21 NET133_22 NET133_23 NET133_24 NET133_25 NET133_26 NET133_27 
+NET133_28 NET133_29 NET133_30 NET133_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 
+BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 
+BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 
+BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 
+BIT_B_29 BIT_B_30 BIT_B_31 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 
+BIT_8 BIT_9 BIT_10 BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 
+BIT_19 BIT_20 BIT_21 BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 
+BIT_30 BIT_31 COL_5 MUX_DEMUX_G17 
XI71 M4_BIT_0 M4_BIT_1 M4_BIT_2 M4_BIT_3 M4_BIT_4 M4_BIT_5 M4_BIT_6 M4_BIT_7 
+M4_BIT_8 M4_BIT_9 M4_BIT_10 M4_BIT_11 M4_BIT_12 M4_BIT_13 M4_BIT_14 M4_BIT_15 
+M4_BIT_16 M4_BIT_17 M4_BIT_18 M4_BIT_19 M4_BIT_20 M4_BIT_21 M4_BIT_22 
+M4_BIT_23 M4_BIT_24 M4_BIT_25 M4_BIT_26 M4_BIT_27 M4_BIT_28 M4_BIT_29 
+M4_BIT_30 M4_BIT_31 M4_BIT_B_0 M4_BIT_B_1 M4_BIT_B_2 M4_BIT_B_3 M4_BIT_B_4 
+M4_BIT_B_5 M4_BIT_B_6 M4_BIT_B_7 M4_BIT_B_8 M4_BIT_B_9 M4_BIT_B_10 M4_BIT_B_11 
+M4_BIT_B_12 M4_BIT_B_13 M4_BIT_B_14 M4_BIT_B_15 M4_BIT_B_16 M4_BIT_B_17 
+M4_BIT_B_18 M4_BIT_B_19 M4_BIT_B_20 M4_BIT_B_21 M4_BIT_B_22 M4_BIT_B_23 
+M4_BIT_B_24 M4_BIT_B_25 M4_BIT_B_26 M4_BIT_B_27 M4_BIT_B_28 M4_BIT_B_29 
+M4_BIT_B_30 M4_BIT_B_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 BIT_B_4 BIT_B_5 
+BIT_B_6 BIT_B_7 BIT_B_8 BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 BIT_B_13 BIT_B_14 
+BIT_B_15 BIT_B_16 BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 BIT_B_21 BIT_B_22 
+BIT_B_23 BIT_B_24 BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 BIT_B_29 BIT_B_30 
+BIT_B_31 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 BIT_8 BIT_9 BIT_10 
+BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 BIT_19 BIT_20 BIT_21 
+BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 BIT_30 BIT_31 COL_4 
+MUX_DEMUX_G17 
XI68 NET199_0 NET199_1 NET199_2 NET199_3 NET199_4 NET199_5 NET199_6 NET199_7 
+NET199_8 NET199_9 NET199_10 NET199_11 NET199_12 NET199_13 NET199_14 NET199_15 
+NET199_16 NET199_17 NET199_18 NET199_19 NET199_20 NET199_21 NET199_22 
+NET199_23 NET199_24 NET199_25 NET199_26 NET199_27 NET199_28 NET199_29 
+NET199_30 NET199_31 NET143_0 NET143_1 NET143_2 NET143_3 NET143_4 NET143_5 
+NET143_6 NET143_7 NET143_8 NET143_9 NET143_10 NET143_11 NET143_12 NET143_13 
+NET143_14 NET143_15 NET143_16 NET143_17 NET143_18 NET143_19 NET143_20 
+NET143_21 NET143_22 NET143_23 NET143_24 NET143_25 NET143_26 NET143_27 
+NET143_28 NET143_29 NET143_30 NET143_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 
+BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 
+BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 
+BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 
+BIT_B_29 BIT_B_30 BIT_B_31 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 
+BIT_8 BIT_9 BIT_10 BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 
+BIT_19 BIT_20 BIT_21 BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 
+BIT_30 BIT_31 COL_1 MUX_DEMUX_G17 
XI73 NET226_0 NET226_1 NET226_2 NET226_3 NET226_4 NET226_5 NET226_6 NET226_7 
+NET226_8 NET226_9 NET226_10 NET226_11 NET226_12 NET226_13 NET226_14 NET226_15 
+NET226_16 NET226_17 NET226_18 NET226_19 NET226_20 NET226_21 NET226_22 
+NET226_23 NET226_24 NET226_25 NET226_26 NET226_27 NET226_28 NET226_29 
+NET226_30 NET226_31 NET148_0 NET148_1 NET148_2 NET148_3 NET148_4 NET148_5 
+NET148_6 NET148_7 NET148_8 NET148_9 NET148_10 NET148_11 NET148_12 NET148_13 
+NET148_14 NET148_15 NET148_16 NET148_17 NET148_18 NET148_19 NET148_20 
+NET148_21 NET148_22 NET148_23 NET148_24 NET148_25 NET148_26 NET148_27 
+NET148_28 NET148_29 NET148_30 NET148_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 
+BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 
+BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 
+BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 
+BIT_B_29 BIT_B_30 BIT_B_31 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 
+BIT_8 BIT_9 BIT_10 BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 
+BIT_19 BIT_20 BIT_21 BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 
+BIT_30 BIT_31 COL_6 MUX_DEMUX_G17 
XI74 NET232_0 NET232_1 NET232_2 NET232_3 NET232_4 NET232_5 NET232_6 NET232_7 
+NET232_8 NET232_9 NET232_10 NET232_11 NET232_12 NET232_13 NET232_14 NET232_15 
+NET232_16 NET232_17 NET232_18 NET232_19 NET232_20 NET232_21 NET232_22 
+NET232_23 NET232_24 NET232_25 NET232_26 NET232_27 NET232_28 NET232_29 
+NET232_30 NET232_31 NET153_0 NET153_1 NET153_2 NET153_3 NET153_4 NET153_5 
+NET153_6 NET153_7 NET153_8 NET153_9 NET153_10 NET153_11 NET153_12 NET153_13 
+NET153_14 NET153_15 NET153_16 NET153_17 NET153_18 NET153_19 NET153_20 
+NET153_21 NET153_22 NET153_23 NET153_24 NET153_25 NET153_26 NET153_27 
+NET153_28 NET153_29 NET153_30 NET153_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 
+BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 
+BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 
+BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 
+BIT_B_29 BIT_B_30 BIT_B_31 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 
+BIT_8 BIT_9 BIT_10 BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 
+BIT_19 BIT_20 BIT_21 BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 
+BIT_30 BIT_31 COL_7 MUX_DEMUX_G17 
XI67 M0_BIT_0 M0_BIT_1 M0_BIT_2 M0_BIT_3 M0_BIT_4 M0_BIT_5 M0_BIT_6 M0_BIT_7 
+M0_BIT_8 M0_BIT_9 M0_BIT_10 M0_BIT_11 M0_BIT_12 M0_BIT_13 M0_BIT_14 M0_BIT_15 
+M0_BIT_16 M0_BIT_17 M0_BIT_18 M0_BIT_19 M0_BIT_20 M0_BIT_21 M0_BIT_22 
+M0_BIT_23 M0_BIT_24 M0_BIT_25 M0_BIT_26 M0_BIT_27 M0_BIT_28 M0_BIT_29 
+M0_BIT_30 M0_BIT_31 M0_BIT_B_0 M0_BIT_B_1 M0_BIT_B_2 M0_BIT_B_3 M0_BIT_B_4 
+M0_BIT_B_5 M0_BIT_B_6 M0_BIT_B_7 M0_BIT_B_8 M0_BIT_B_9 M0_BIT_B_10 M0_BIT_B_11 
+M0_BIT_B_12 M0_BIT_B_13 M0_BIT_B_14 M0_BIT_B_15 M0_BIT_B_16 M0_BIT_B_17 
+M0_BIT_B_18 M0_BIT_B_19 M0_BIT_B_20 M0_BIT_B_21 M0_BIT_B_22 M0_BIT_B_23 
+M0_BIT_B_24 M0_BIT_B_25 M0_BIT_B_26 M0_BIT_B_27 M0_BIT_B_28 M0_BIT_B_29 
+M0_BIT_B_30 M0_BIT_B_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 BIT_B_4 BIT_B_5 
+BIT_B_6 BIT_B_7 BIT_B_8 BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 BIT_B_13 BIT_B_14 
+BIT_B_15 BIT_B_16 BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 BIT_B_21 BIT_B_22 
+BIT_B_23 BIT_B_24 BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 BIT_B_29 BIT_B_30 
+BIT_B_31 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 BIT_8 BIT_9 BIT_10 
+BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 BIT_19 BIT_20 BIT_21 
+BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 BIT_30 BIT_31 COL_0 
+MUX_DEMUX_G17 
XI69 NET205_0 NET205_1 NET205_2 NET205_3 NET205_4 NET205_5 NET205_6 NET205_7 
+NET205_8 NET205_9 NET205_10 NET205_11 NET205_12 NET205_13 NET205_14 NET205_15 
+NET205_16 NET205_17 NET205_18 NET205_19 NET205_20 NET205_21 NET205_22 
+NET205_23 NET205_24 NET205_25 NET205_26 NET205_27 NET205_28 NET205_29 
+NET205_30 NET205_31 NET163_0 NET163_1 NET163_2 NET163_3 NET163_4 NET163_5 
+NET163_6 NET163_7 NET163_8 NET163_9 NET163_10 NET163_11 NET163_12 NET163_13 
+NET163_14 NET163_15 NET163_16 NET163_17 NET163_18 NET163_19 NET163_20 
+NET163_21 NET163_22 NET163_23 NET163_24 NET163_25 NET163_26 NET163_27 
+NET163_28 NET163_29 NET163_30 NET163_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 
+BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 
+BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 
+BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 
+BIT_B_29 BIT_B_30 BIT_B_31 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 
+BIT_8 BIT_9 BIT_10 BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 
+BIT_19 BIT_20 BIT_21 BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 
+BIT_30 BIT_31 COL_2 MUX_DEMUX_G17 
XI70 NET214_0 NET214_1 NET214_2 NET214_3 NET214_4 NET214_5 NET214_6 NET214_7 
+NET214_8 NET214_9 NET214_10 NET214_11 NET214_12 NET214_13 NET214_14 NET214_15 
+NET214_16 NET214_17 NET214_18 NET214_19 NET214_20 NET214_21 NET214_22 
+NET214_23 NET214_24 NET214_25 NET214_26 NET214_27 NET214_28 NET214_29 
+NET214_30 NET214_31 NET168_0 NET168_1 NET168_2 NET168_3 NET168_4 NET168_5 
+NET168_6 NET168_7 NET168_8 NET168_9 NET168_10 NET168_11 NET168_12 NET168_13 
+NET168_14 NET168_15 NET168_16 NET168_17 NET168_18 NET168_19 NET168_20 
+NET168_21 NET168_22 NET168_23 NET168_24 NET168_25 NET168_26 NET168_27 
+NET168_28 NET168_29 NET168_30 NET168_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 
+BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 
+BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 
+BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 
+BIT_B_29 BIT_B_30 BIT_B_31 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 
+BIT_8 BIT_9 BIT_10 BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 
+BIT_19 BIT_20 BIT_21 BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 
+BIT_30 BIT_31 COL_3 MUX_DEMUX_G17 
XI63 ADDRESS_A_7 ADDRESS_A_8 ADDRESS_A_9 ADDRESS_B_7 ADDRESS_B_8 ADDRESS_B_9 
+COL_0 COL_1 COL_2 COL_3 COL_4 COL_5 COL_6 COL_7 COL_DEC_G18 
XI47 WL_A_0 WL_A_1 WL_A_2 WL_A_3 WL_A_4 WL_A_5 WL_A_6 WL_A_7 WL_A_8 WL_A_9 
+WL_A_10 WL_A_11 WL_A_12 WL_A_13 WL_A_14 WL_A_15 WL_A_16 WL_A_17 WL_A_18 
+WL_A_19 WL_A_20 WL_A_21 WL_A_22 WL_A_23 WL_A_24 WL_A_25 WL_A_26 WL_A_27 
+WL_A_28 WL_A_29 WL_A_30 WL_A_31 WL_A_32 WL_A_33 WL_A_34 WL_A_35 WL_A_36 
+WL_A_37 WL_A_38 WL_A_39 WL_A_40 WL_A_41 WL_A_42 WL_A_43 WL_A_44 WL_A_45 
+WL_A_46 WL_A_47 WL_A_48 WL_A_49 WL_A_50 WL_A_51 WL_A_52 WL_A_53 WL_A_54 
+WL_A_55 WL_A_56 WL_A_57 WL_A_58 WL_A_59 WL_A_60 WL_A_61 WL_A_62 WL_A_63 WL_B_0 
+WL_B_1 WL_B_2 WL_B_3 WL_B_4 WL_B_5 WL_B_6 WL_B_7 WL_B_8 WL_B_9 WL_B_10 WL_B_11 
+WL_B_12 WL_B_13 WL_B_14 WL_B_15 WL_B_16 WL_B_17 WL_B_18 WL_B_19 WL_B_20 
+WL_B_21 WL_B_22 WL_B_23 WL_B_24 WL_B_25 WL_B_26 WL_B_27 WL_B_28 WL_B_29 
+WL_B_30 WL_B_31 WL_B_32 WL_B_33 WL_B_34 WL_B_35 WL_B_36 WL_B_37 WL_B_38 
+WL_B_39 WL_B_40 WL_B_41 WL_B_42 WL_B_43 WL_B_44 WL_B_45 WL_B_46 WL_B_47 
+WL_B_48 WL_B_49 WL_B_50 WL_B_51 WL_B_52 WL_B_53 WL_B_54 WL_B_55 WL_B_56 
+WL_B_57 WL_B_58 WL_B_59 WL_B_60 WL_B_61 WL_B_62 WL_B_63 WORD_EN_REAL 
+CONTROL_G19 
XI48 WL_A_64 WL_A_65 WL_A_66 WL_A_67 WL_A_68 WL_A_69 WL_A_70 WL_A_71 WL_A_72 
+WL_A_73 WL_A_74 WL_A_75 WL_A_76 WL_A_77 WL_A_78 WL_A_79 WL_A_80 WL_A_81 
+WL_A_82 WL_A_83 WL_A_84 WL_A_85 WL_A_86 WL_A_87 WL_A_88 WL_A_89 WL_A_90 
+WL_A_91 WL_A_92 WL_A_93 WL_A_94 WL_A_95 WL_A_96 WL_A_97 WL_A_98 WL_A_99 
+WL_A_100 WL_A_101 WL_A_102 WL_A_103 WL_A_104 WL_A_105 WL_A_106 WL_A_107 
+WL_A_108 WL_A_109 WL_A_110 WL_A_111 WL_A_112 WL_A_113 WL_A_114 WL_A_115 
+WL_A_116 WL_A_117 WL_A_118 WL_A_119 WL_A_120 WL_A_121 WL_A_122 WL_A_123 
+WL_A_124 WL_A_125 WL_A_126 WL_A_127 WL_B_64 WL_B_65 WL_B_66 WL_B_67 WL_B_68 
+WL_B_69 WL_B_70 WL_B_71 WL_B_72 WL_B_73 WL_B_74 WL_B_75 WL_B_76 WL_B_77 
+WL_B_78 WL_B_79 WL_B_80 WL_B_81 WL_B_82 WL_B_83 WL_B_84 WL_B_85 WL_B_86 
+WL_B_87 WL_B_88 WL_B_89 WL_B_90 WL_B_91 WL_B_92 WL_B_93 WL_B_94 WL_B_95 
+WL_B_96 WL_B_97 WL_B_98 WL_B_99 WL_B_100 WL_B_101 WL_B_102 WL_B_103 WL_B_104 
+WL_B_105 WL_B_106 WL_B_107 WL_B_108 WL_B_109 WL_B_110 WL_B_111 WL_B_112 
+WL_B_113 WL_B_114 WL_B_115 WL_B_116 WL_B_117 WL_B_118 WL_B_119 WL_B_120 
+WL_B_121 WL_B_122 WL_B_123 WL_B_124 WL_B_125 WL_B_126 WL_B_127 WORD_EN_REAL 
+CONTROL_G19 
XI46 ADDRESS_A_0 ADDRESS_A_1 ADDRESS_A_2 ADDRESS_A_3 ADDRESS_A_4 ADDRESS_A_5 
+ADDRESS_A_6 ADDRESS_BUF_0 ADDRESS_BUF_1 ADDRESS_BUF_2 ADDRESS_BUF_3 
+ADDRESS_BUF_4 ADDRESS_BUF_5 ADDRESS_BUF_6 ADDRESS_B_0 ADDRESS_B_1 ADDRESS_B_2 
+ADDRESS_B_3 ADDRESS_B_4 ADDRESS_B_5 ADDRESS_B_6 PATH1INVS7_G20 
XI45 CLK ADDRESS_0 ADDRESS_1 ADDRESS_2 ADDRESS_3 ADDRESS_4 ADDRESS_5 ADDRESS_6 
+ADDRESS_7 ADDRESS_8 ADDRESS_9 NET0104_0 NET0104_1 NET0104_2 NET0104_3 
+NET0104_4 NET0104_5 NET0104_6 NET0105_0 NET0105_1 NET0105_2 REG10_G21 
XI43 WL_B_0 WL_B_1 WL_B_2 WL_B_3 WL_B_4 WL_B_5 WL_B_6 WL_B_7 WL_B_8 WL_B_9 
+WL_B_10 WL_B_11 WL_B_12 WL_B_13 WL_B_14 WL_B_15 WL_B_16 WL_B_17 WL_B_18 
+WL_B_19 WL_B_20 WL_B_21 WL_B_22 WL_B_23 WL_B_24 WL_B_25 WL_B_26 WL_B_27 
+WL_B_28 WL_B_29 WL_B_30 WL_B_31 WL_B_32 WL_B_33 WL_B_34 WL_B_35 WL_B_36 
+WL_B_37 WL_B_38 WL_B_39 WL_B_40 WL_B_41 WL_B_42 WL_B_43 WL_B_44 WL_B_45 
+WL_B_46 WL_B_47 WL_B_48 WL_B_49 WL_B_50 WL_B_51 WL_B_52 WL_B_53 WL_B_54 
+WL_B_55 WL_B_56 WL_B_57 WL_B_58 WL_B_59 WL_B_60 WL_B_61 WL_B_62 WL_B_63 WL_0 
+WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 
+WL_15 WL_16 WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 
+WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 
+WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 
+WL_54 WL_55 WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 SUB1 
XI44 WL_B_64 WL_B_65 WL_B_66 WL_B_67 WL_B_68 WL_B_69 WL_B_70 WL_B_71 WL_B_72 
+WL_B_73 WL_B_74 WL_B_75 WL_B_76 WL_B_77 WL_B_78 WL_B_79 WL_B_80 WL_B_81 
+WL_B_82 WL_B_83 WL_B_84 WL_B_85 WL_B_86 WL_B_87 WL_B_88 WL_B_89 WL_B_90 
+WL_B_91 WL_B_92 WL_B_93 WL_B_94 WL_B_95 WL_B_96 WL_B_97 WL_B_98 WL_B_99 
+WL_B_100 WL_B_101 WL_B_102 WL_B_103 WL_B_104 WL_B_105 WL_B_106 WL_B_107 
+WL_B_108 WL_B_109 WL_B_110 WL_B_111 WL_B_112 WL_B_113 WL_B_114 WL_B_115 
+WL_B_116 WL_B_117 WL_B_118 WL_B_119 WL_B_120 WL_B_121 WL_B_122 WL_B_123 
+WL_B_124 WL_B_125 WL_B_126 WL_B_127 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 
+WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 
+WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 
+WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 
+WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118 
+WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 SUB1 
XI42 WL_A_0 WL_A_1 WL_A_2 WL_A_3 WL_A_4 WL_A_5 WL_A_6 WL_A_7 WL_A_8 WL_A_9 
+WL_A_10 WL_A_11 WL_A_12 WL_A_13 WL_A_14 WL_A_15 WL_A_16 WL_A_17 WL_A_18 
+WL_A_19 WL_A_20 WL_A_21 WL_A_22 WL_A_23 WL_A_24 WL_A_25 WL_A_26 WL_A_27 
+WL_A_28 WL_A_29 WL_A_30 WL_A_31 WL_A_32 WL_A_33 WL_A_34 WL_A_35 WL_A_36 
+WL_A_37 WL_A_38 WL_A_39 WL_A_40 WL_A_41 WL_A_42 WL_A_43 WL_A_44 WL_A_45 
+WL_A_46 WL_A_47 WL_A_48 WL_A_49 WL_A_50 WL_A_51 WL_A_52 WL_A_53 WL_A_54 
+WL_A_55 WL_A_56 WL_A_57 WL_A_58 WL_A_59 WL_A_60 WL_A_61 WL_A_62 WL_A_63 
+WL_A_64 WL_A_65 WL_A_66 WL_A_67 WL_A_68 WL_A_69 WL_A_70 WL_A_71 WL_A_72 
+WL_A_73 WL_A_74 WL_A_75 WL_A_76 WL_A_77 WL_A_78 WL_A_79 WL_A_80 WL_A_81 
+WL_A_82 WL_A_83 WL_A_84 WL_A_85 WL_A_86 WL_A_87 WL_A_88 WL_A_89 WL_A_90 
+WL_A_91 WL_A_92 WL_A_93 WL_A_94 WL_A_95 WL_A_96 WL_A_97 WL_A_98 WL_A_99 
+WL_A_100 WL_A_101 WL_A_102 WL_A_103 WL_A_104 WL_A_105 WL_A_106 WL_A_107 
+WL_A_108 WL_A_109 WL_A_110 WL_A_111 WL_A_112 WL_A_113 WL_A_114 WL_A_115 
+WL_A_116 WL_A_117 WL_A_118 WL_A_119 WL_A_120 WL_A_121 WL_A_122 WL_A_123 
+WL_A_124 WL_A_125 WL_A_126 WL_A_127 ADDRESS_BUF_0 ADDRESS_BUF_1 ADDRESS_BUF_2 
+ADDRESS_BUF_3 ADDRESS_BUF_4 ADDRESS_BUF_5 ADDRESS_BUF_6 ADDRESS_B_0 
+ADDRESS_B_1 ADDRESS_B_2 ADDRESS_B_3 ADDRESS_B_4 ADDRESS_B_5 ADDRESS_B_6 
+RDEC7TO128_G22 
XI49 NET199_0 NET199_1 NET199_2 NET199_3 NET199_4 NET199_5 NET199_6 NET199_7 
+NET199_8 NET199_9 NET199_10 NET199_11 NET199_12 NET199_13 NET199_14 NET199_15 
+NET199_16 NET199_17 NET199_18 NET199_19 NET199_20 NET199_21 NET199_22 
+NET199_23 NET199_24 NET199_25 NET199_26 NET199_27 NET199_28 NET199_29 
+NET199_30 NET199_31 NET143_0 NET143_1 NET143_2 NET143_3 NET143_4 NET143_5 
+NET143_6 NET143_7 NET143_8 NET143_9 NET143_10 NET143_11 NET143_12 NET143_13 
+NET143_14 NET143_15 NET143_16 NET143_17 NET143_18 NET143_19 NET143_20 
+NET143_21 NET143_22 NET143_23 NET143_24 NET143_25 NET143_26 NET143_27 
+NET143_28 NET143_29 NET143_30 NET143_31 WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 
+WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18 WL_19 
+WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 
+WL_33 WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 
+WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58 
+WL_59 WL_60 WL_61 WL_62 WL_63 SUB2 
XI50 NET199_0 NET199_1 NET199_2 NET199_3 NET199_4 NET199_5 NET199_6 NET199_7 
+NET199_8 NET199_9 NET199_10 NET199_11 NET199_12 NET199_13 NET199_14 NET199_15 
+NET199_16 NET199_17 NET199_18 NET199_19 NET199_20 NET199_21 NET199_22 
+NET199_23 NET199_24 NET199_25 NET199_26 NET199_27 NET199_28 NET199_29 
+NET199_30 NET199_31 NET143_0 NET143_1 NET143_2 NET143_3 NET143_4 NET143_5 
+NET143_6 NET143_7 NET143_8 NET143_9 NET143_10 NET143_11 NET143_12 NET143_13 
+NET143_14 NET143_15 NET143_16 NET143_17 NET143_18 NET143_19 NET143_20 
+NET143_21 NET143_22 NET143_23 NET143_24 NET143_25 NET143_26 NET143_27 
+NET143_28 NET143_29 NET143_30 NET143_31 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 
+WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 
+WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 
+WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 
+WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 
+WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 SUB2 
XI51 NET205_0 NET205_1 NET205_2 NET205_3 NET205_4 NET205_5 NET205_6 NET205_7 
+NET205_8 NET205_9 NET205_10 NET205_11 NET205_12 NET205_13 NET205_14 NET205_15 
+NET205_16 NET205_17 NET205_18 NET205_19 NET205_20 NET205_21 NET205_22 
+NET205_23 NET205_24 NET205_25 NET205_26 NET205_27 NET205_28 NET205_29 
+NET205_30 NET205_31 NET163_0 NET163_1 NET163_2 NET163_3 NET163_4 NET163_5 
+NET163_6 NET163_7 NET163_8 NET163_9 NET163_10 NET163_11 NET163_12 NET163_13 
+NET163_14 NET163_15 NET163_16 NET163_17 NET163_18 NET163_19 NET163_20 
+NET163_21 NET163_22 NET163_23 NET163_24 NET163_25 NET163_26 NET163_27 
+NET163_28 NET163_29 NET163_30 NET163_31 WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 
+WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18 WL_19 
+WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 
+WL_33 WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 
+WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58 
+WL_59 WL_60 WL_61 WL_62 WL_63 SUB2 
XI52 NET205_0 NET205_1 NET205_2 NET205_3 NET205_4 NET205_5 NET205_6 NET205_7 
+NET205_8 NET205_9 NET205_10 NET205_11 NET205_12 NET205_13 NET205_14 NET205_15 
+NET205_16 NET205_17 NET205_18 NET205_19 NET205_20 NET205_21 NET205_22 
+NET205_23 NET205_24 NET205_25 NET205_26 NET205_27 NET205_28 NET205_29 
+NET205_30 NET205_31 NET163_0 NET163_1 NET163_2 NET163_3 NET163_4 NET163_5 
+NET163_6 NET163_7 NET163_8 NET163_9 NET163_10 NET163_11 NET163_12 NET163_13 
+NET163_14 NET163_15 NET163_16 NET163_17 NET163_18 NET163_19 NET163_20 
+NET163_21 NET163_22 NET163_23 NET163_24 NET163_25 NET163_26 NET163_27 
+NET163_28 NET163_29 NET163_30 NET163_31 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 
+WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 
+WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 
+WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 
+WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 
+WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 SUB2 
XSRAM4BOT M4_BIT_0 M4_BIT_1 M4_BIT_2 M4_BIT_3 M4_BIT_4 M4_BIT_5 M4_BIT_6 
+M4_BIT_7 M4_BIT_8 M4_BIT_9 M4_BIT_10 M4_BIT_11 M4_BIT_12 M4_BIT_13 M4_BIT_14 
+M4_BIT_15 M4_BIT_16 M4_BIT_17 M4_BIT_18 M4_BIT_19 M4_BIT_20 M4_BIT_21 
+M4_BIT_22 M4_BIT_23 M4_BIT_24 M4_BIT_25 M4_BIT_26 M4_BIT_27 M4_BIT_28 
+M4_BIT_29 M4_BIT_30 M4_BIT_31 M4_BIT_B_0 M4_BIT_B_1 M4_BIT_B_2 M4_BIT_B_3 
+M4_BIT_B_4 M4_BIT_B_5 M4_BIT_B_6 M4_BIT_B_7 M4_BIT_B_8 M4_BIT_B_9 M4_BIT_B_10 
+M4_BIT_B_11 M4_BIT_B_12 M4_BIT_B_13 M4_BIT_B_14 M4_BIT_B_15 M4_BIT_B_16 
+M4_BIT_B_17 M4_BIT_B_18 M4_BIT_B_19 M4_BIT_B_20 M4_BIT_B_21 M4_BIT_B_22 
+M4_BIT_B_23 M4_BIT_B_24 M4_BIT_B_25 M4_BIT_B_26 M4_BIT_B_27 M4_BIT_B_28 
+M4_BIT_B_29 M4_BIT_B_30 M4_BIT_B_31 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 
+WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 
+WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 
+WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 
+WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118 
+WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 SUB2 
XI58 NET220_0 NET220_1 NET220_2 NET220_3 NET220_4 NET220_5 NET220_6 NET220_7 
+NET220_8 NET220_9 NET220_10 NET220_11 NET220_12 NET220_13 NET220_14 NET220_15 
+NET220_16 NET220_17 NET220_18 NET220_19 NET220_20 NET220_21 NET220_22 
+NET220_23 NET220_24 NET220_25 NET220_26 NET220_27 NET220_28 NET220_29 
+NET220_30 NET220_31 NET133_0 NET133_1 NET133_2 NET133_3 NET133_4 NET133_5 
+NET133_6 NET133_7 NET133_8 NET133_9 NET133_10 NET133_11 NET133_12 NET133_13 
+NET133_14 NET133_15 NET133_16 NET133_17 NET133_18 NET133_19 NET133_20 
+NET133_21 NET133_22 NET133_23 NET133_24 NET133_25 NET133_26 NET133_27 
+NET133_28 NET133_29 NET133_30 NET133_31 WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 
+WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18 WL_19 
+WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 
+WL_33 WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 
+WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58 
+WL_59 WL_60 WL_61 WL_62 WL_63 SUB2 
XI53 NET214_0 NET214_1 NET214_2 NET214_3 NET214_4 NET214_5 NET214_6 NET214_7 
+NET214_8 NET214_9 NET214_10 NET214_11 NET214_12 NET214_13 NET214_14 NET214_15 
+NET214_16 NET214_17 NET214_18 NET214_19 NET214_20 NET214_21 NET214_22 
+NET214_23 NET214_24 NET214_25 NET214_26 NET214_27 NET214_28 NET214_29 
+NET214_30 NET214_31 NET168_0 NET168_1 NET168_2 NET168_3 NET168_4 NET168_5 
+NET168_6 NET168_7 NET168_8 NET168_9 NET168_10 NET168_11 NET168_12 NET168_13 
+NET168_14 NET168_15 NET168_16 NET168_17 NET168_18 NET168_19 NET168_20 
+NET168_21 NET168_22 NET168_23 NET168_24 NET168_25 NET168_26 NET168_27 
+NET168_28 NET168_29 NET168_30 NET168_31 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 
+WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 
+WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 
+WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 
+WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 
+WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 SUB2 
XI54 NET214_0 NET214_1 NET214_2 NET214_3 NET214_4 NET214_5 NET214_6 NET214_7 
+NET214_8 NET214_9 NET214_10 NET214_11 NET214_12 NET214_13 NET214_14 NET214_15 
+NET214_16 NET214_17 NET214_18 NET214_19 NET214_20 NET214_21 NET214_22 
+NET214_23 NET214_24 NET214_25 NET214_26 NET214_27 NET214_28 NET214_29 
+NET214_30 NET214_31 NET168_0 NET168_1 NET168_2 NET168_3 NET168_4 NET168_5 
+NET168_6 NET168_7 NET168_8 NET168_9 NET168_10 NET168_11 NET168_12 NET168_13 
+NET168_14 NET168_15 NET168_16 NET168_17 NET168_18 NET168_19 NET168_20 
+NET168_21 NET168_22 NET168_23 NET168_24 NET168_25 NET168_26 NET168_27 
+NET168_28 NET168_29 NET168_30 NET168_31 WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 
+WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18 WL_19 
+WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 
+WL_33 WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 
+WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58 
+WL_59 WL_60 WL_61 WL_62 WL_63 SUB2 
XI57 NET220_0 NET220_1 NET220_2 NET220_3 NET220_4 NET220_5 NET220_6 NET220_7 
+NET220_8 NET220_9 NET220_10 NET220_11 NET220_12 NET220_13 NET220_14 NET220_15 
+NET220_16 NET220_17 NET220_18 NET220_19 NET220_20 NET220_21 NET220_22 
+NET220_23 NET220_24 NET220_25 NET220_26 NET220_27 NET220_28 NET220_29 
+NET220_30 NET220_31 NET133_0 NET133_1 NET133_2 NET133_3 NET133_4 NET133_5 
+NET133_6 NET133_7 NET133_8 NET133_9 NET133_10 NET133_11 NET133_12 NET133_13 
+NET133_14 NET133_15 NET133_16 NET133_17 NET133_18 NET133_19 NET133_20 
+NET133_21 NET133_22 NET133_23 NET133_24 NET133_25 NET133_26 NET133_27 
+NET133_28 NET133_29 NET133_30 NET133_31 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 
+WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 
+WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 
+WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 
+WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 
+WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 SUB2 
XSRAM0BOT M0_BIT_0 M0_BIT_1 M0_BIT_2 M0_BIT_3 M0_BIT_4 M0_BIT_5 M0_BIT_6 
+M0_BIT_7 M0_BIT_8 M0_BIT_9 M0_BIT_10 M0_BIT_11 M0_BIT_12 M0_BIT_13 M0_BIT_14 
+M0_BIT_15 M0_BIT_16 M0_BIT_17 M0_BIT_18 M0_BIT_19 M0_BIT_20 M0_BIT_21 
+M0_BIT_22 M0_BIT_23 M0_BIT_24 M0_BIT_25 M0_BIT_26 M0_BIT_27 M0_BIT_28 
+M0_BIT_29 M0_BIT_30 M0_BIT_31 M0_BIT_B_0 M0_BIT_B_1 M0_BIT_B_2 M0_BIT_B_3 
+M0_BIT_B_4 M0_BIT_B_5 M0_BIT_B_6 M0_BIT_B_7 M0_BIT_B_8 M0_BIT_B_9 M0_BIT_B_10 
+M0_BIT_B_11 M0_BIT_B_12 M0_BIT_B_13 M0_BIT_B_14 M0_BIT_B_15 M0_BIT_B_16 
+M0_BIT_B_17 M0_BIT_B_18 M0_BIT_B_19 M0_BIT_B_20 M0_BIT_B_21 M0_BIT_B_22 
+M0_BIT_B_23 M0_BIT_B_24 M0_BIT_B_25 M0_BIT_B_26 M0_BIT_B_27 M0_BIT_B_28 
+M0_BIT_B_29 M0_BIT_B_30 M0_BIT_B_31 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 WL_70 
+WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 WL_83 
+WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 WL_96 
+WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 WL_107 
+WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 WL_118 
+WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 SUB2 
XI59 NET226_0 NET226_1 NET226_2 NET226_3 NET226_4 NET226_5 NET226_6 NET226_7 
+NET226_8 NET226_9 NET226_10 NET226_11 NET226_12 NET226_13 NET226_14 NET226_15 
+NET226_16 NET226_17 NET226_18 NET226_19 NET226_20 NET226_21 NET226_22 
+NET226_23 NET226_24 NET226_25 NET226_26 NET226_27 NET226_28 NET226_29 
+NET226_30 NET226_31 NET148_0 NET148_1 NET148_2 NET148_3 NET148_4 NET148_5 
+NET148_6 NET148_7 NET148_8 NET148_9 NET148_10 NET148_11 NET148_12 NET148_13 
+NET148_14 NET148_15 NET148_16 NET148_17 NET148_18 NET148_19 NET148_20 
+NET148_21 NET148_22 NET148_23 NET148_24 NET148_25 NET148_26 NET148_27 
+NET148_28 NET148_29 NET148_30 NET148_31 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 
+WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 
+WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 
+WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 
+WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 
+WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 SUB2 
XI60 NET226_0 NET226_1 NET226_2 NET226_3 NET226_4 NET226_5 NET226_6 NET226_7 
+NET226_8 NET226_9 NET226_10 NET226_11 NET226_12 NET226_13 NET226_14 NET226_15 
+NET226_16 NET226_17 NET226_18 NET226_19 NET226_20 NET226_21 NET226_22 
+NET226_23 NET226_24 NET226_25 NET226_26 NET226_27 NET226_28 NET226_29 
+NET226_30 NET226_31 NET148_0 NET148_1 NET148_2 NET148_3 NET148_4 NET148_5 
+NET148_6 NET148_7 NET148_8 NET148_9 NET148_10 NET148_11 NET148_12 NET148_13 
+NET148_14 NET148_15 NET148_16 NET148_17 NET148_18 NET148_19 NET148_20 
+NET148_21 NET148_22 NET148_23 NET148_24 NET148_25 NET148_26 NET148_27 
+NET148_28 NET148_29 NET148_30 NET148_31 WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 
+WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18 WL_19 
+WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 
+WL_33 WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 
+WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58 
+WL_59 WL_60 WL_61 WL_62 WL_63 SUB2 
XI61 NET232_0 NET232_1 NET232_2 NET232_3 NET232_4 NET232_5 NET232_6 NET232_7 
+NET232_8 NET232_9 NET232_10 NET232_11 NET232_12 NET232_13 NET232_14 NET232_15 
+NET232_16 NET232_17 NET232_18 NET232_19 NET232_20 NET232_21 NET232_22 
+NET232_23 NET232_24 NET232_25 NET232_26 NET232_27 NET232_28 NET232_29 
+NET232_30 NET232_31 NET153_0 NET153_1 NET153_2 NET153_3 NET153_4 NET153_5 
+NET153_6 NET153_7 NET153_8 NET153_9 NET153_10 NET153_11 NET153_12 NET153_13 
+NET153_14 NET153_15 NET153_16 NET153_17 NET153_18 NET153_19 NET153_20 
+NET153_21 NET153_22 NET153_23 NET153_24 NET153_25 NET153_26 NET153_27 
+NET153_28 NET153_29 NET153_30 NET153_31 WL_64 WL_65 WL_66 WL_67 WL_68 WL_69 
+WL_70 WL_71 WL_72 WL_73 WL_74 WL_75 WL_76 WL_77 WL_78 WL_79 WL_80 WL_81 WL_82 
+WL_83 WL_84 WL_85 WL_86 WL_87 WL_88 WL_89 WL_90 WL_91 WL_92 WL_93 WL_94 WL_95 
+WL_96 WL_97 WL_98 WL_99 WL_100 WL_101 WL_102 WL_103 WL_104 WL_105 WL_106 
+WL_107 WL_108 WL_109 WL_110 WL_111 WL_112 WL_113 WL_114 WL_115 WL_116 WL_117 
+WL_118 WL_119 WL_120 WL_121 WL_122 WL_123 WL_124 WL_125 WL_126 WL_127 SUB2 
XI62 NET232_0 NET232_1 NET232_2 NET232_3 NET232_4 NET232_5 NET232_6 NET232_7 
+NET232_8 NET232_9 NET232_10 NET232_11 NET232_12 NET232_13 NET232_14 NET232_15 
+NET232_16 NET232_17 NET232_18 NET232_19 NET232_20 NET232_21 NET232_22 
+NET232_23 NET232_24 NET232_25 NET232_26 NET232_27 NET232_28 NET232_29 
+NET232_30 NET232_31 NET153_0 NET153_1 NET153_2 NET153_3 NET153_4 NET153_5 
+NET153_6 NET153_7 NET153_8 NET153_9 NET153_10 NET153_11 NET153_12 NET153_13 
+NET153_14 NET153_15 NET153_16 NET153_17 NET153_18 NET153_19 NET153_20 
+NET153_21 NET153_22 NET153_23 NET153_24 NET153_25 NET153_26 NET153_27 
+NET153_28 NET153_29 NET153_30 NET153_31 WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 
+WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18 WL_19 
+WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 
+WL_33 WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 
+WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58 
+WL_59 WL_60 WL_61 WL_62 WL_63 SUB2 
XSRAM4TOP M4_BIT_0 M4_BIT_1 M4_BIT_2 M4_BIT_3 M4_BIT_4 M4_BIT_5 M4_BIT_6 
+M4_BIT_7 M4_BIT_8 M4_BIT_9 M4_BIT_10 M4_BIT_11 M4_BIT_12 M4_BIT_13 M4_BIT_14 
+M4_BIT_15 M4_BIT_16 M4_BIT_17 M4_BIT_18 M4_BIT_19 M4_BIT_20 M4_BIT_21 
+M4_BIT_22 M4_BIT_23 M4_BIT_24 M4_BIT_25 M4_BIT_26 M4_BIT_27 M4_BIT_28 
+M4_BIT_29 M4_BIT_30 M4_BIT_31 M4_BIT_B_0 M4_BIT_B_1 M4_BIT_B_2 M4_BIT_B_3 
+M4_BIT_B_4 M4_BIT_B_5 M4_BIT_B_6 M4_BIT_B_7 M4_BIT_B_8 M4_BIT_B_9 M4_BIT_B_10 
+M4_BIT_B_11 M4_BIT_B_12 M4_BIT_B_13 M4_BIT_B_14 M4_BIT_B_15 M4_BIT_B_16 
+M4_BIT_B_17 M4_BIT_B_18 M4_BIT_B_19 M4_BIT_B_20 M4_BIT_B_21 M4_BIT_B_22 
+M4_BIT_B_23 M4_BIT_B_24 M4_BIT_B_25 M4_BIT_B_26 M4_BIT_B_27 M4_BIT_B_28 
+M4_BIT_B_29 M4_BIT_B_30 M4_BIT_B_31 WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 
+WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18 WL_19 WL_20 
+WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 
+WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 
+WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58 WL_59 
+WL_60 WL_61 WL_62 WL_63 SUB2 
XSRAM0TOP M0_BIT_0 M0_BIT_1 M0_BIT_2 M0_BIT_3 M0_BIT_4 M0_BIT_5 M0_BIT_6 
+M0_BIT_7 M0_BIT_8 M0_BIT_9 M0_BIT_10 M0_BIT_11 M0_BIT_12 M0_BIT_13 M0_BIT_14 
+M0_BIT_15 M0_BIT_16 M0_BIT_17 M0_BIT_18 M0_BIT_19 M0_BIT_20 M0_BIT_21 
+M0_BIT_22 M0_BIT_23 M0_BIT_24 M0_BIT_25 M0_BIT_26 M0_BIT_27 M0_BIT_28 
+M0_BIT_29 M0_BIT_30 M0_BIT_31 M0_BIT_B_0 M0_BIT_B_1 M0_BIT_B_2 M0_BIT_B_3 
+M0_BIT_B_4 M0_BIT_B_5 M0_BIT_B_6 M0_BIT_B_7 M0_BIT_B_8 M0_BIT_B_9 M0_BIT_B_10 
+M0_BIT_B_11 M0_BIT_B_12 M0_BIT_B_13 M0_BIT_B_14 M0_BIT_B_15 M0_BIT_B_16 
+M0_BIT_B_17 M0_BIT_B_18 M0_BIT_B_19 M0_BIT_B_20 M0_BIT_B_21 M0_BIT_B_22 
+M0_BIT_B_23 M0_BIT_B_24 M0_BIT_B_25 M0_BIT_B_26 M0_BIT_B_27 M0_BIT_B_28 
+M0_BIT_B_29 M0_BIT_B_30 M0_BIT_B_31 WL_0 WL_1 WL_2 WL_3 WL_4 WL_5 WL_6 WL_7 
+WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 WL_17 WL_18 WL_19 WL_20 
+WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 WL_30 WL_31 WL_32 WL_33 
+WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 WL_43 WL_44 WL_45 WL_46 
+WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 WL_56 WL_57 WL_58 WL_59 
+WL_60 WL_61 WL_62 WL_63 SUB2 
XI64 ADDRESS_A_7 ADDRESS_B_7 INV_5 
XI65 ADDRESS_A_8 ADDRESS_B_8 INV_5 
XI66 ADDRESS_A_9 ADDRESS_B_9 INV_5 
XI12 NET112_0 NET112_1 NET112_2 NET112_3 NET112_4 NET112_5 NET112_6 NET112_7 
+NET112_8 NET112_9 NET112_10 NET112_11 NET112_12 NET112_13 NET112_14 NET112_15 
+NET112_16 NET112_17 NET112_18 NET112_19 NET112_20 NET112_21 NET112_22 
+NET112_23 NET112_24 NET112_25 NET112_26 NET112_27 NET112_28 NET112_29 
+NET112_30 NET112_31 NET254_0 NET254_1 NET254_2 NET254_3 NET254_4 NET254_5 
+NET254_6 NET254_7 NET254_8 NET254_9 NET254_10 NET254_11 NET254_12 NET254_13 
+NET254_14 NET254_15 NET254_16 NET254_17 NET254_18 NET254_19 NET254_20 
+NET254_21 NET254_22 NET254_23 NET254_24 NET254_25 NET254_26 NET254_27 
+NET254_28 NET254_29 NET254_30 NET254_31 INV32_G23 
XI16 CLK NET257_0 NET257_1 NET257_2 NET257_3 NET257_4 NET257_5 NET257_6 
+NET257_7 NET257_8 NET257_9 NET257_10 NET257_11 NET257_12 NET257_13 NET257_14 
+NET257_15 NET257_16 NET257_17 NET257_18 NET257_19 NET257_20 NET257_21 
+NET257_22 NET257_23 NET257_24 NET257_25 NET257_26 NET257_27 NET257_28 
+NET257_29 NET257_30 NET257_31 DATA_OUT_B_0 DATA_OUT_B_1 DATA_OUT_B_2 
+DATA_OUT_B_3 DATA_OUT_B_4 DATA_OUT_B_5 DATA_OUT_B_6 DATA_OUT_B_7 DATA_OUT_B_8 
+DATA_OUT_B_9 DATA_OUT_B_10 DATA_OUT_B_11 DATA_OUT_B_12 DATA_OUT_B_13 
+DATA_OUT_B_14 DATA_OUT_B_15 DATA_OUT_B_16 DATA_OUT_B_17 DATA_OUT_B_18 
+DATA_OUT_B_19 DATA_OUT_B_20 DATA_OUT_B_21 DATA_OUT_B_22 DATA_OUT_B_23 
+DATA_OUT_B_24 DATA_OUT_B_25 DATA_OUT_B_26 DATA_OUT_B_27 DATA_OUT_B_28 
+DATA_OUT_B_29 DATA_OUT_B_30 DATA_OUT_B_31 REG32_G24 
XI15 CLK NET260_0 NET260_1 NET260_2 NET260_3 NET260_4 NET260_5 NET260_6 
+NET260_7 NET260_8 NET260_9 NET260_10 NET260_11 NET260_12 NET260_13 NET260_14 
+NET260_15 NET260_16 NET260_17 NET260_18 NET260_19 NET260_20 NET260_21 
+NET260_22 NET260_23 NET260_24 NET260_25 NET260_26 NET260_27 NET260_28 
+NET260_29 NET260_30 NET260_31 DATA_OUT_0 DATA_OUT_1 DATA_OUT_2 DATA_OUT_3 
+DATA_OUT_4 DATA_OUT_5 DATA_OUT_6 DATA_OUT_7 DATA_OUT_8 DATA_OUT_9 DATA_OUT_10 
+DATA_OUT_11 DATA_OUT_12 DATA_OUT_13 DATA_OUT_14 DATA_OUT_15 DATA_OUT_16 
+DATA_OUT_17 DATA_OUT_18 DATA_OUT_19 DATA_OUT_20 DATA_OUT_21 DATA_OUT_22 
+DATA_OUT_23 DATA_OUT_24 DATA_OUT_25 DATA_OUT_26 DATA_OUT_27 DATA_OUT_28 
+DATA_OUT_29 DATA_OUT_30 DATA_OUT_31 REG32_G24 
XI6 CLK DATA_IN_0 DATA_IN_1 DATA_IN_2 DATA_IN_3 DATA_IN_4 DATA_IN_5 DATA_IN_6 
+DATA_IN_7 DATA_IN_8 DATA_IN_9 DATA_IN_10 DATA_IN_11 DATA_IN_12 DATA_IN_13 
+DATA_IN_14 DATA_IN_15 DATA_IN_16 DATA_IN_17 DATA_IN_18 DATA_IN_19 DATA_IN_20 
+DATA_IN_21 DATA_IN_22 DATA_IN_23 DATA_IN_24 DATA_IN_25 DATA_IN_26 DATA_IN_27 
+DATA_IN_28 DATA_IN_29 DATA_IN_30 DATA_IN_31 NET262_0 NET262_1 NET262_2 
+NET262_3 NET262_4 NET262_5 NET262_6 NET262_7 NET262_8 NET262_9 NET262_10 
+NET262_11 NET262_12 NET262_13 NET262_14 NET262_15 NET262_16 NET262_17 
+NET262_18 NET262_19 NET262_20 NET262_21 NET262_22 NET262_23 NET262_24 
+NET262_25 NET262_26 NET262_27 NET262_28 NET262_29 NET262_30 NET262_31 
+REG32_G24 
XI3 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 BIT_8 BIT_9 BIT_10 BIT_11 
+BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 BIT_19 BIT_20 BIT_21 BIT_22 
+BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 BIT_30 BIT_31 BIT_0 BIT_1 
+BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 BIT_8 BIT_9 BIT_10 BIT_11 BIT_12 BIT_13 
+BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 BIT_19 BIT_20 BIT_21 BIT_22 BIT_23 BIT_24 
+BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 BIT_30 BIT_31 BIT_B_0 BIT_B_1 BIT_B_2 
+BIT_B_3 BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 BIT_B_9 BIT_B_10 BIT_B_11 
+BIT_B_12 BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 BIT_B_17 BIT_B_18 BIT_B_19 
+BIT_B_20 BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 BIT_B_25 BIT_B_26 BIT_B_27 
+BIT_B_28 BIT_B_29 BIT_B_30 BIT_B_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 BIT_B_4 
+BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 BIT_B_13 
+BIT_B_14 BIT_B_15 BIT_B_16 BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 BIT_B_21 
+BIT_B_22 BIT_B_23 BIT_B_24 BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 BIT_B_29 
+BIT_B_30 BIT_B_31 NET112_0 NET112_1 NET112_2 NET112_3 NET112_4 NET112_5 
+NET112_6 NET112_7 NET112_8 NET112_9 NET112_10 NET112_11 NET112_12 NET112_13 
+NET112_14 NET112_15 NET112_16 NET112_17 NET112_18 NET112_19 NET112_20 
+NET112_21 NET112_22 NET112_23 NET112_24 NET112_25 NET112_26 NET112_27 
+NET112_28 NET112_29 NET112_30 NET112_31 NET254_0 NET254_1 NET254_2 NET254_3 
+NET254_4 NET254_5 NET254_6 NET254_7 NET254_8 NET254_9 NET254_10 NET254_11 
+NET254_12 NET254_13 NET254_14 NET254_15 NET254_16 NET254_17 NET254_18 
+NET254_19 NET254_20 NET254_21 NET254_22 NET254_23 NET254_24 NET254_25 
+NET254_26 NET254_27 NET254_28 NET254_29 NET254_30 NET254_31 PRE_REAL 
+WRITE_EN_REAL WRITE_CELL32_G25 
XSENSEAMP BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 BIT_8 BIT_9 BIT_10 
+BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 BIT_19 BIT_20 BIT_21 
+BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 BIT_30 BIT_31 BIT_B_0 
+BIT_B_1 BIT_B_2 BIT_B_3 BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 BIT_B_9 
+BIT_B_10 BIT_B_11 BIT_B_12 BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 BIT_B_17 
+BIT_B_18 BIT_B_19 BIT_B_20 BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 BIT_B_25 
+BIT_B_26 BIT_B_27 BIT_B_28 BIT_B_29 BIT_B_30 BIT_B_31 NET116_0 NET116_1 
+NET116_2 NET116_3 NET116_4 NET116_5 NET116_6 NET116_7 NET116_8 NET116_9 
+NET116_10 NET116_11 NET116_12 NET116_13 NET116_14 NET116_15 NET116_16 
+NET116_17 NET116_18 NET116_19 NET116_20 NET116_21 NET116_22 NET116_23 
+NET116_24 NET116_25 NET116_26 NET116_27 NET116_28 NET116_29 NET116_30 
+NET116_31 OUT_B_PRE_FF_0 OUT_B_PRE_FF_1 OUT_B_PRE_FF_2 OUT_B_PRE_FF_3 
+OUT_B_PRE_FF_4 OUT_B_PRE_FF_5 OUT_B_PRE_FF_6 OUT_B_PRE_FF_7 OUT_B_PRE_FF_8 
+OUT_B_PRE_FF_9 OUT_B_PRE_FF_10 OUT_B_PRE_FF_11 OUT_B_PRE_FF_12 OUT_B_PRE_FF_13 
+OUT_B_PRE_FF_14 OUT_B_PRE_FF_15 OUT_B_PRE_FF_16 OUT_B_PRE_FF_17 
+OUT_B_PRE_FF_18 OUT_B_PRE_FF_19 OUT_B_PRE_FF_20 OUT_B_PRE_FF_21 
+OUT_B_PRE_FF_22 OUT_B_PRE_FF_23 OUT_B_PRE_FF_24 OUT_B_PRE_FF_25 
+OUT_B_PRE_FF_26 OUT_B_PRE_FF_27 OUT_B_PRE_FF_28 OUT_B_PRE_FF_29 
+OUT_B_PRE_FF_30 OUT_B_PRE_FF_31 READ_EN_REAL SAMP_CELL32_G26 
   
* FILE NAME: SRAM2_TL_PI_MODEL32_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL32.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN<0> = IN_0
*                   IN<1> = IN_1
*                   IN<2> = IN_2
*                   IN<3> = IN_3
*                   IN<4> = IN_4
*                   IN<5> = IN_5
*                   IN<6> = IN_6
*                   IN<7> = IN_7
*                   IN<8> = IN_8
*                   IN<9> = IN_9
*                   IN<10> = IN_10
*                   IN<11> = IN_11
*                   IN<12> = IN_12
*                   IN<13> = IN_13
*                   IN<14> = IN_14
*                   IN<15> = IN_15
*                   IN<16> = IN_16
*                   IN<17> = IN_17
*                   IN<18> = IN_18
*                   IN<19> = IN_19
*                   IN<20> = IN_20
*                   IN<21> = IN_21
*                   IN<22> = IN_22
*                   IN<23> = IN_23
*                   IN<24> = IN_24
*                   IN<25> = IN_25
*                   IN<26> = IN_26
*                   IN<27> = IN_27
*                   IN<28> = IN_28
*                   IN<29> = IN_29
*                   IN<30> = IN_30
*                   IN<31> = IN_31
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
*                   OUT<3> = OUT_3
*                   OUT<4> = OUT_4
*                   OUT<5> = OUT_5
*                   OUT<6> = OUT_6
*                   OUT<7> = OUT_7
*                   OUT<8> = OUT_8
*                   OUT<9> = OUT_9
*                   OUT<10> = OUT_10
*                   OUT<11> = OUT_11
*                   OUT<12> = OUT_12
*                   OUT<13> = OUT_13
*                   OUT<14> = OUT_14
*                   OUT<15> = OUT_15
*                   OUT<16> = OUT_16
*                   OUT<17> = OUT_17
*                   OUT<18> = OUT_18
*                   OUT<19> = OUT_19
*                   OUT<20> = OUT_20
*                   OUT<21> = OUT_21
*                   OUT<22> = OUT_22
*                   OUT<23> = OUT_23
*                   OUT<24> = OUT_24
*                   OUT<25> = OUT_25
*                   OUT<26> = OUT_26
*                   OUT<27> = OUT_27
*                   OUT<28> = OUT_28
*                   OUT<29> = OUT_29
*                   OUT<30> = OUT_30
*                   OUT<31> = OUT_31
.SUBCKT TL_PI_MODEL32_3 IN_0 IN_1 IN_2 IN_3 IN_4 IN_5 IN_6 IN_7 IN_8 IN_9 
+IN_10 IN_11 IN_12 IN_13 IN_14 IN_15 IN_16 IN_17 IN_18 IN_19 IN_20 IN_21 IN_22 
+IN_23 IN_24 IN_25 IN_26 IN_27 IN_28 IN_29 IN_30 IN_31 OUT_0 OUT_1 OUT_2 OUT_3 
+OUT_4 OUT_5 OUT_6 OUT_7 OUT_8 OUT_9 OUT_10 OUT_11 OUT_12 OUT_13 OUT_14 OUT_15 
+OUT_16 OUT_17 OUT_18 OUT_19 OUT_20 OUT_21 OUT_22 OUT_23 OUT_24 OUT_25 OUT_26 
+OUT_27 OUT_28 OUT_29 OUT_30 OUT_31 
XI31 IN_31 OUT_31 TL_PI_MODEL_1 
XI30 IN_30 OUT_30 TL_PI_MODEL_1 
XI29 IN_29 OUT_29 TL_PI_MODEL_1 
XI28 IN_28 OUT_28 TL_PI_MODEL_1 
XI27 IN_27 OUT_27 TL_PI_MODEL_1 
XI26 IN_26 OUT_26 TL_PI_MODEL_1 
XI25 IN_25 OUT_25 TL_PI_MODEL_1 
XI24 IN_24 OUT_24 TL_PI_MODEL_1 
XI23 IN_23 OUT_23 TL_PI_MODEL_1 
XI22 IN_22 OUT_22 TL_PI_MODEL_1 
XI21 IN_21 OUT_21 TL_PI_MODEL_1 
XI20 IN_20 OUT_20 TL_PI_MODEL_1 
XI19 IN_19 OUT_19 TL_PI_MODEL_1 
XI18 IN_18 OUT_18 TL_PI_MODEL_1 
XI17 IN_17 OUT_17 TL_PI_MODEL_1 
XI16 IN_16 OUT_16 TL_PI_MODEL_1 
XI15 IN_15 OUT_15 TL_PI_MODEL_1 
XI14 IN_14 OUT_14 TL_PI_MODEL_1 
XI13 IN_13 OUT_13 TL_PI_MODEL_1 
XI12 IN_12 OUT_12 TL_PI_MODEL_1 
XI11 IN_11 OUT_11 TL_PI_MODEL_1 
XI10 IN_10 OUT_10 TL_PI_MODEL_1 
XI9 IN_9 OUT_9 TL_PI_MODEL_1 
XI8 IN_8 OUT_8 TL_PI_MODEL_1 
XI7 IN_7 OUT_7 TL_PI_MODEL_1 
XI6 IN_6 OUT_6 TL_PI_MODEL_1 
XI5 IN_5 OUT_5 TL_PI_MODEL_1 
XI4 IN_4 OUT_4 TL_PI_MODEL_1 
XI3 IN_3 OUT_3 TL_PI_MODEL_1 
XI2 IN_2 OUT_2 TL_PI_MODEL_1 
XI1 IN_1 OUT_1 TL_PI_MODEL_1 
XI0 IN_0 OUT_0 TL_PI_MODEL_1 
   
   
* FILE NAME: SRAM2_TL_PI_MODEL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:31 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT TL_PI_MODEL_1 IN OUT 
C0 IN 0  ((33E-15)) M=1.0 
C1 OUT 0  ((33E-15)) M=1.0 
R0 IN OUT  ((115.2)) M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL32_3 
* FILE NAME: SRAM2_TL_PI_MODEL32_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL32.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN<0> = IN_0
*                   IN<1> = IN_1
*                   IN<2> = IN_2
*                   IN<3> = IN_3
*                   IN<4> = IN_4
*                   IN<5> = IN_5
*                   IN<6> = IN_6
*                   IN<7> = IN_7
*                   IN<8> = IN_8
*                   IN<9> = IN_9
*                   IN<10> = IN_10
*                   IN<11> = IN_11
*                   IN<12> = IN_12
*                   IN<13> = IN_13
*                   IN<14> = IN_14
*                   IN<15> = IN_15
*                   IN<16> = IN_16
*                   IN<17> = IN_17
*                   IN<18> = IN_18
*                   IN<19> = IN_19
*                   IN<20> = IN_20
*                   IN<21> = IN_21
*                   IN<22> = IN_22
*                   IN<23> = IN_23
*                   IN<24> = IN_24
*                   IN<25> = IN_25
*                   IN<26> = IN_26
*                   IN<27> = IN_27
*                   IN<28> = IN_28
*                   IN<29> = IN_29
*                   IN<30> = IN_30
*                   IN<31> = IN_31
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
*                   OUT<3> = OUT_3
*                   OUT<4> = OUT_4
*                   OUT<5> = OUT_5
*                   OUT<6> = OUT_6
*                   OUT<7> = OUT_7
*                   OUT<8> = OUT_8
*                   OUT<9> = OUT_9
*                   OUT<10> = OUT_10
*                   OUT<11> = OUT_11
*                   OUT<12> = OUT_12
*                   OUT<13> = OUT_13
*                   OUT<14> = OUT_14
*                   OUT<15> = OUT_15
*                   OUT<16> = OUT_16
*                   OUT<17> = OUT_17
*                   OUT<18> = OUT_18
*                   OUT<19> = OUT_19
*                   OUT<20> = OUT_20
*                   OUT<21> = OUT_21
*                   OUT<22> = OUT_22
*                   OUT<23> = OUT_23
*                   OUT<24> = OUT_24
*                   OUT<25> = OUT_25
*                   OUT<26> = OUT_26
*                   OUT<27> = OUT_27
*                   OUT<28> = OUT_28
*                   OUT<29> = OUT_29
*                   OUT<30> = OUT_30
*                   OUT<31> = OUT_31
.SUBCKT TL_PI_MODEL32_4 IN_0 IN_1 IN_2 IN_3 IN_4 IN_5 IN_6 IN_7 IN_8 IN_9 
+IN_10 IN_11 IN_12 IN_13 IN_14 IN_15 IN_16 IN_17 IN_18 IN_19 IN_20 IN_21 IN_22 
+IN_23 IN_24 IN_25 IN_26 IN_27 IN_28 IN_29 IN_30 IN_31 OUT_0 OUT_1 OUT_2 OUT_3 
+OUT_4 OUT_5 OUT_6 OUT_7 OUT_8 OUT_9 OUT_10 OUT_11 OUT_12 OUT_13 OUT_14 OUT_15 
+OUT_16 OUT_17 OUT_18 OUT_19 OUT_20 OUT_21 OUT_22 OUT_23 OUT_24 OUT_25 OUT_26 
+OUT_27 OUT_28 OUT_29 OUT_30 OUT_31 
XI31 IN_31 OUT_31 TL_PI_MODEL_1 
XI30 IN_30 OUT_30 TL_PI_MODEL_1 
XI29 IN_29 OUT_29 TL_PI_MODEL_1 
XI28 IN_28 OUT_28 TL_PI_MODEL_1 
XI27 IN_27 OUT_27 TL_PI_MODEL_1 
XI26 IN_26 OUT_26 TL_PI_MODEL_1 
XI25 IN_25 OUT_25 TL_PI_MODEL_1 
XI24 IN_24 OUT_24 TL_PI_MODEL_1 
XI23 IN_23 OUT_23 TL_PI_MODEL_1 
XI22 IN_22 OUT_22 TL_PI_MODEL_1 
XI21 IN_21 OUT_21 TL_PI_MODEL_1 
XI20 IN_20 OUT_20 TL_PI_MODEL_1 
XI19 IN_19 OUT_19 TL_PI_MODEL_1 
XI18 IN_18 OUT_18 TL_PI_MODEL_1 
XI17 IN_17 OUT_17 TL_PI_MODEL_1 
XI16 IN_16 OUT_16 TL_PI_MODEL_1 
XI15 IN_15 OUT_15 TL_PI_MODEL_1 
XI14 IN_14 OUT_14 TL_PI_MODEL_1 
XI13 IN_13 OUT_13 TL_PI_MODEL_1 
XI12 IN_12 OUT_12 TL_PI_MODEL_1 
XI11 IN_11 OUT_11 TL_PI_MODEL_1 
XI10 IN_10 OUT_10 TL_PI_MODEL_1 
XI9 IN_9 OUT_9 TL_PI_MODEL_1 
XI8 IN_8 OUT_8 TL_PI_MODEL_1 
XI7 IN_7 OUT_7 TL_PI_MODEL_1 
XI6 IN_6 OUT_6 TL_PI_MODEL_1 
XI5 IN_5 OUT_5 TL_PI_MODEL_1 
XI4 IN_4 OUT_4 TL_PI_MODEL_1 
XI3 IN_3 OUT_3 TL_PI_MODEL_1 
XI2 IN_2 OUT_2 TL_PI_MODEL_1 
XI1 IN_1 OUT_1 TL_PI_MODEL_1 
XI0 IN_0 OUT_0 TL_PI_MODEL_1 
   
   
* FILE NAME: SRAM2_TL_PI_MODEL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:31 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT TL_PI_MODEL_1 IN OUT 
C0 IN 0  ((33.5E-15)) M=1.0 
C1 OUT 0  ((33.5E-15)) M=1.0 
R0 IN OUT  ((153.6)) M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL32_4 
* FILE NAME: SRAM2_TL_PI_MODEL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:31 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT TL_PI_MODEL_2 IN OUT 
C0 IN 0  (34.6E-15) M=1.0 
C1 OUT 0  (34.6E-15) M=1.0 
R0 IN OUT  (230.4) M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL_2 
* FILE NAME: SRAM2_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_5 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(18E-6) AD=+9.00000000E-12 
+AS=+9.00000000E-12 PD=+3.70000000E-05 PS=+3.70000000E-05 NRD=+2.77777778E-02 
+NRS=+2.77777778E-02 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(6E-6) AD=+3.00000000E-12 AS=+3.00000000E-12 
+PD=+1.30000000E-05 PS=+1.30000000E-05 NRD=+8.33333333E-02 NRS=+8.33333333E-02 
+M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_5 
* FILE NAME: SRAM2_TL_PI_MODEL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:31 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT TL_PI_MODEL_1 IN OUT 
C0 IN 0  (33E-15) M=1.0 
C1 OUT 0  (33E-15) M=1.0 
R0 IN OUT  (128.0) M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL_1 
   
   
   
* FILE NAME: SRAM2_DUMMY_ROW_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: DUMMY_ROW.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:33 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   PRE_REAL = PRE_REAL
*                   READ_EN_REAL = READ_EN_REAL
*                   WORD_EN_REAL = WORD_EN_REAL
*                   WRITE_EN = WRITE_EN
.SUBCKT DUMMY_ROW_G15 CLK PRE_REAL READ_EN_REAL WORD_EN_REAL WRITE_EN 
M0 DUM_BIT DUM_WL VDD! VDD!  PFET  L=200E-9 W=800E-9 AD=+4.00000000E-13 
+AS=+4.00000000E-13 PD=+2.60000000E-06 PS=+2.60000000E-06 NRD=+6.25000000E-01 
+NRS=+6.25000000E-01 M=1.0 
XI195 DELAY_B CLK NET035 NAND2_1 
XI169 NET051 CLK_B NET038 NAND2_1 
XI86 NET040 DELAY_B NET055 NAND2_2 
XI203 NET035 NET043 INV_3 
XI197 NET043 PRE_REAL INV_3 
XI201 NET044 WORD_EN_REAL INV_3 
XI200 DELAY NET044 INV_4 
XI177 WRITE_EN NET051 INV_4 
XI202 NET055 READ_EN_REAL INV_3 
XI196 NET038 NET040 INV_4 
XI199 DELAY_B DELAY INV_4 
XI198 DUM_BIT DELAY_B INV_4 
XI156 CLK CLK_B INV_5 
XI150 CLK_B DUM_WL TL_PI_MODEL_6 
XI139 DUM_BIT NET42 DUM_WL NET40 DUM_SRAM_CELL_G2 
XI193 DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT NET0111_0 NET0111_1 NET0111_2 
+NET0111_3 NET0111_4 NET0111_5 NET0111_6 NET0111_7 NET0111_8 NET0111_9 
+NET0111_10 NET0111_11 NET0111_12 NET0111_13 NET0111_14 NET0111_15 NET0111_16 
+NET0111_17 NET0111_18 NET0111_19 NET0111_20 NET0111_21 NET0111_22 NET0111_23 
+NET0111_24 NET0111_25 NET0111_26 NET0111_27 NET0111_28 NET0111_29 NET0111_30 
+NET0111_31 0 SRAM_CELL32_G3 
XI192 DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT NET0114_0 NET0114_1 NET0114_2 
+NET0114_3 NET0114_4 NET0114_5 NET0114_6 NET0114_7 NET0114_8 NET0114_9 
+NET0114_10 NET0114_11 NET0114_12 NET0114_13 NET0114_14 NET0114_15 NET0114_16 
+NET0114_17 NET0114_18 NET0114_19 NET0114_20 NET0114_21 NET0114_22 NET0114_23 
+NET0114_24 NET0114_25 NET0114_26 NET0114_27 NET0114_28 NET0114_29 NET0114_30 
+NET0114_31 0 SRAM_CELL32_G3 
XI191 DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT NET0117_0 NET0117_1 NET0117_2 
+NET0117_3 NET0117_4 NET0117_5 NET0117_6 NET0117_7 NET0117_8 NET0117_9 
+NET0117_10 NET0117_11 NET0117_12 NET0117_13 NET0117_14 NET0117_15 NET0117_16 
+NET0117_17 NET0117_18 NET0117_19 NET0117_20 NET0117_21 NET0117_22 NET0117_23 
+NET0117_24 NET0117_25 NET0117_26 NET0117_27 NET0117_28 NET0117_29 NET0117_30 
+NET0117_31 0 SRAM_CELL32_G3 
XI190 DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT 
+DUM_BIT DUM_BIT DUM_BIT DUM_BIT DUM_BIT NET0120_0 NET0120_1 NET0120_2 
+NET0120_3 NET0120_4 NET0120_5 NET0120_6 NET0120_7 NET0120_8 NET0120_9 
+NET0120_10 NET0120_11 NET0120_12 NET0120_13 NET0120_14 NET0120_15 NET0120_16 
+NET0120_17 NET0120_18 NET0120_19 NET0120_20 NET0120_21 NET0120_22 NET0120_23 
+NET0120_24 NET0120_25 NET0120_26 NET0120_27 NET0120_28 NET0120_29 NET0120_30 
+NET0120_31 0 SRAM_CELL32_G3 
XI9 NET80_0 NET80_1 NET80_2 NET80_3 NET80_4 NET80_5 NET80_6 NET80_7 NET80_8 
+NET80_9 NET80_10 NET80_11 NET80_12 NET80_13 NET80_14 NET80_15 NET80_16 
+NET80_17 NET80_18 NET80_19 NET80_20 NET80_21 NET80_22 NET80_23 NET80_24 
+NET80_25 NET80_26 NET80_27 NET80_28 NET80_29 NET80_30 NET80_31 NET81_0 NET81_1 
+NET81_2 NET81_3 NET81_4 NET81_5 NET81_6 NET81_7 NET81_8 NET81_9 NET81_10 
+NET81_11 NET81_12 NET81_13 NET81_14 NET81_15 NET81_16 NET81_17 NET81_18 
+NET81_19 NET81_20 NET81_21 NET81_22 NET81_23 NET81_24 NET81_25 NET81_26 
+NET81_27 NET81_28 NET81_29 NET81_30 NET81_31 DUM_WL SRAM_CELL32_G3 
XI8 NET83_0 NET83_1 NET83_2 NET83_3 NET83_4 NET83_5 NET83_6 NET83_7 NET83_8 
+NET83_9 NET83_10 NET83_11 NET83_12 NET83_13 NET83_14 NET83_15 NET83_16 
+NET83_17 NET83_18 NET83_19 NET83_20 NET83_21 NET83_22 NET83_23 NET83_24 
+NET83_25 NET83_26 NET83_27 NET83_28 NET83_29 NET83_30 NET83_31 NET84_0 NET84_1 
+NET84_2 NET84_3 NET84_4 NET84_5 NET84_6 NET84_7 NET84_8 NET84_9 NET84_10 
+NET84_11 NET84_12 NET84_13 NET84_14 NET84_15 NET84_16 NET84_17 NET84_18 
+NET84_19 NET84_20 NET84_21 NET84_22 NET84_23 NET84_24 NET84_25 NET84_26 
+NET84_27 NET84_28 NET84_29 NET84_30 NET84_31 DUM_WL SRAM_CELL32_G3 
XI7 NET86_0 NET86_1 NET86_2 NET86_3 NET86_4 NET86_5 NET86_6 NET86_7 NET86_8 
+NET86_9 NET86_10 NET86_11 NET86_12 NET86_13 NET86_14 NET86_15 NET86_16 
+NET86_17 NET86_18 NET86_19 NET86_20 NET86_21 NET86_22 NET86_23 NET86_24 
+NET86_25 NET86_26 NET86_27 NET86_28 NET86_29 NET86_30 NET86_31 NET87_0 NET87_1 
+NET87_2 NET87_3 NET87_4 NET87_5 NET87_6 NET87_7 NET87_8 NET87_9 NET87_10 
+NET87_11 NET87_12 NET87_13 NET87_14 NET87_15 NET87_16 NET87_17 NET87_18 
+NET87_19 NET87_20 NET87_21 NET87_22 NET87_23 NET87_24 NET87_25 NET87_26 
+NET87_27 NET87_28 NET87_29 NET87_30 NET87_31 DUM_WL SRAM_CELL32_G3 
XI6 NET89_0 NET89_1 NET89_2 NET89_3 NET89_4 NET89_5 NET89_6 NET89_7 NET89_8 
+NET89_9 NET89_10 NET89_11 NET89_12 NET89_13 NET89_14 NET89_15 NET89_16 
+NET89_17 NET89_18 NET89_19 NET89_20 NET89_21 NET89_22 NET89_23 NET89_24 
+NET89_25 NET89_26 NET89_27 NET89_28 NET89_29 NET89_30 NET89_31 NET90_0 NET90_1 
+NET90_2 NET90_3 NET90_4 NET90_5 NET90_6 NET90_7 NET90_8 NET90_9 NET90_10 
+NET90_11 NET90_12 NET90_13 NET90_14 NET90_15 NET90_16 NET90_17 NET90_18 
+NET90_19 NET90_20 NET90_21 NET90_22 NET90_23 NET90_24 NET90_25 NET90_26 
+NET90_27 NET90_28 NET90_29 NET90_30 NET90_31 DUM_WL SRAM_CELL32_G3 
XI4 NET92_0 NET92_1 NET92_2 NET92_3 NET92_4 NET92_5 NET92_6 NET92_7 NET92_8 
+NET92_9 NET92_10 NET92_11 NET92_12 NET92_13 NET92_14 NET92_15 NET92_16 
+NET92_17 NET92_18 NET92_19 NET92_20 NET92_21 NET92_22 NET92_23 NET92_24 
+NET92_25 NET92_26 NET92_27 NET92_28 NET92_29 NET92_30 NET92_31 NET93_0 NET93_1 
+NET93_2 NET93_3 NET93_4 NET93_5 NET93_6 NET93_7 NET93_8 NET93_9 NET93_10 
+NET93_11 NET93_12 NET93_13 NET93_14 NET93_15 NET93_16 NET93_17 NET93_18 
+NET93_19 NET93_20 NET93_21 NET93_22 NET93_23 NET93_24 NET93_25 NET93_26 
+NET93_27 NET93_28 NET93_29 NET93_30 NET93_31 DUM_WL SRAM_CELL32_G3 
   
   
* FILE NAME: SRAM2_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_5 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(48.1E-6) AD=+2.40500000E-11 
+AS=+2.40500000E-11 PD=+9.72000000E-05 PS=+9.72000000E-05 NRD=+1.03950104E-02 
+NRS=+1.03950104E-02 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(16E-6) AD=+8.00000000E-12 AS=+8.00000000E-12 
+PD=+3.30000000E-05 PS=+3.30000000E-05 NRD=+3.12500000E-02 NRS=+3.12500000E-02 
+M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_5 
* FILE NAME: SRAM2_NAND2_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: NAND2.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   OUT = OUT
.SUBCKT NAND2_1 A B OUT 
M3 OUT B VDD! VDD!  PFET  L=200E-9 W=(27E-6) AD=+1.35000000E-11 
+AS=+1.35000000E-11 PD=+5.50000000E-05 PS=+5.50000000E-05 NRD=+1.85185185E-02 
+NRS=+1.85185185E-02 M=1.0 
M2 OUT A VDD! VDD!  PFET  L=200E-9 W=(27E-6) AD=+1.35000000E-11 
+AS=+1.35000000E-11 PD=+5.50000000E-05 PS=+5.50000000E-05 NRD=+1.85185185E-02 
+NRS=+1.85185185E-02 M=1.0 
M1 OUT A NET15 0  NFET  L=200E-9 W=(18E-6) AD=+9.00000000E-12 
+AS=+9.00000000E-12 PD=+3.70000000E-05 PS=+3.70000000E-05 NRD=+2.77777778E-02 
+NRS=+2.77777778E-02 M=1.0 
M0 NET15 B 0 0  NFET  L=200E-9 W=(18E-6) AD=+9.00000000E-12 AS=+9.00000000E-12 
+PD=+3.70000000E-05 PS=+3.70000000E-05 NRD=+2.77777778E-02 NRS=+2.77777778E-02 
+M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NAND2_1 
* FILE NAME: SRAM2_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_3 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(270E-6) AD=+1.35000000E-10 
+AS=+1.35000000E-10 PD=+5.41000000E-04 PS=+5.41000000E-04 NRD=+1.85185185E-03 
+NRS=+1.85185185E-03 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(90E-6) AD=+4.50000000E-11 AS=+4.50000000E-11 
+PD=+1.81000000E-04 PS=+1.81000000E-04 NRD=+5.55555556E-03 NRS=+5.55555556E-03 
+M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_3 
* FILE NAME: SRAM2_TL_PI_MODEL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:31 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT TL_PI_MODEL_6 IN OUT 
C0 IN 0  (291E-15) M=1.0 
C1 OUT 0  (291E-15) M=1.0 
R0 IN OUT  (204.8) M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL_6 
* FILE NAME: SRAM2_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_4 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(27E-6) AD=+1.35000000E-11 
+AS=+1.35000000E-11 PD=+5.50000000E-05 PS=+5.50000000E-05 NRD=+1.85185185E-02 
+NRS=+1.85185185E-02 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(9E-6) AD=+4.50000000E-12 AS=+4.50000000E-12 
+PD=+1.90000000E-05 PS=+1.90000000E-05 NRD=+5.55555556E-02 NRS=+5.55555556E-02 
+M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_4 
* FILE NAME: SRAM2_NAND2_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: NAND2.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   OUT = OUT
.SUBCKT NAND2_2 A B OUT 
M3 OUT B VDD! VDD!  PFET  L=200E-9 W=(102E-6) AD=+5.10000000E-11 
+AS=+5.10000000E-11 PD=+2.05000000E-04 PS=+2.05000000E-04 NRD=+4.90196078E-03 
+NRS=+4.90196078E-03 M=1.0 
M2 OUT A VDD! VDD!  PFET  L=200E-9 W=(102E-6) AD=+5.10000000E-11 
+AS=+5.10000000E-11 PD=+2.05000000E-04 PS=+2.05000000E-04 NRD=+4.90196078E-03 
+NRS=+4.90196078E-03 M=1.0 
M1 OUT A NET15 0  NFET  L=200E-9 W=(68E-6) AD=+3.40000000E-11 
+AS=+3.40000000E-11 PD=+1.37000000E-04 PS=+1.37000000E-04 NRD=+7.35294118E-03 
+NRS=+7.35294118E-03 M=1.0 
M0 NET15 B 0 0  NFET  L=200E-9 W=(68E-6) AD=+3.40000000E-11 AS=+3.40000000E-11 
+PD=+1.37000000E-04 PS=+1.37000000E-04 NRD=+7.35294118E-03 NRS=+7.35294118E-03 
+M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NAND2_2 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS DUMMY_ROW_G15 
* FILE NAME: SRAM2_SRAM_CELL32_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SRAM_CELL32.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: BIT<0> = BIT_0
*                   BIT<1> = BIT_1
*                   BIT<2> = BIT_2
*                   BIT<3> = BIT_3
*                   BIT<4> = BIT_4
*                   BIT<5> = BIT_5
*                   BIT<6> = BIT_6
*                   BIT<7> = BIT_7
*                   BIT<8> = BIT_8
*                   BIT<9> = BIT_9
*                   BIT<10> = BIT_10
*                   BIT<11> = BIT_11
*                   BIT<12> = BIT_12
*                   BIT<13> = BIT_13
*                   BIT<14> = BIT_14
*                   BIT<15> = BIT_15
*                   BIT<16> = BIT_16
*                   BIT<17> = BIT_17
*                   BIT<18> = BIT_18
*                   BIT<19> = BIT_19
*                   BIT<20> = BIT_20
*                   BIT<21> = BIT_21
*                   BIT<22> = BIT_22
*                   BIT<23> = BIT_23
*                   BIT<24> = BIT_24
*                   BIT<25> = BIT_25
*                   BIT<26> = BIT_26
*                   BIT<27> = BIT_27
*                   BIT<28> = BIT_28
*                   BIT<29> = BIT_29
*                   BIT<30> = BIT_30
*                   BIT<31> = BIT_31
*                   BIT_B<0> = BIT_B_0
*                   BIT_B<1> = BIT_B_1
*                   BIT_B<2> = BIT_B_2
*                   BIT_B<3> = BIT_B_3
*                   BIT_B<4> = BIT_B_4
*                   BIT_B<5> = BIT_B_5
*                   BIT_B<6> = BIT_B_6
*                   BIT_B<7> = BIT_B_7
*                   BIT_B<8> = BIT_B_8
*                   BIT_B<9> = BIT_B_9
*                   BIT_B<10> = BIT_B_10
*                   BIT_B<11> = BIT_B_11
*                   BIT_B<12> = BIT_B_12
*                   BIT_B<13> = BIT_B_13
*                   BIT_B<14> = BIT_B_14
*                   BIT_B<15> = BIT_B_15
*                   BIT_B<16> = BIT_B_16
*                   BIT_B<17> = BIT_B_17
*                   BIT_B<18> = BIT_B_18
*                   BIT_B<19> = BIT_B_19
*                   BIT_B<20> = BIT_B_20
*                   BIT_B<21> = BIT_B_21
*                   BIT_B<22> = BIT_B_22
*                   BIT_B<23> = BIT_B_23
*                   BIT_B<24> = BIT_B_24
*                   BIT_B<25> = BIT_B_25
*                   BIT_B<26> = BIT_B_26
*                   BIT_B<27> = BIT_B_27
*                   BIT_B<28> = BIT_B_28
*                   BIT_B<29> = BIT_B_29
*                   BIT_B<30> = BIT_B_30
*                   BIT_B<31> = BIT_B_31
*                   WL = WL
.SUBCKT SRAM_CELL32_G3 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 BIT_8 
+BIT_9 BIT_10 BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 BIT_19 
+BIT_20 BIT_21 BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 BIT_30 
+BIT_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 
+BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 
+BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 
+BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 BIT_B_29 BIT_B_30 BIT_B_31 WL 
XI32 BIT_31 NET101 NET100 WL BIT_B_31 SRAM_CELL_G1 
XI31 BIT_30 NET106 NET105 WL BIT_B_30 SRAM_CELL_G1 
XI30 BIT_29 NET111 NET110 WL BIT_B_29 SRAM_CELL_G1 
XI29 BIT_28 NET116 NET115 WL BIT_B_28 SRAM_CELL_G1 
XI28 BIT_27 NET121 NET120 WL BIT_B_27 SRAM_CELL_G1 
XI27 BIT_26 NET126 NET125 WL BIT_B_26 SRAM_CELL_G1 
XI26 BIT_25 NET131 NET130 WL BIT_B_25 SRAM_CELL_G1 
XI25 BIT_24 NET136 NET135 WL BIT_B_24 SRAM_CELL_G1 
XI24 BIT_23 NET141 NET140 WL BIT_B_23 SRAM_CELL_G1 
XI23 BIT_22 NET146 NET145 WL BIT_B_22 SRAM_CELL_G1 
XI22 BIT_21 NET151 NET150 WL BIT_B_21 SRAM_CELL_G1 
XI21 BIT_20 NET156 NET155 WL BIT_B_20 SRAM_CELL_G1 
XI20 BIT_19 NET161 NET160 WL BIT_B_19 SRAM_CELL_G1 
XI19 BIT_18 NET166 NET165 WL BIT_B_18 SRAM_CELL_G1 
XI18 BIT_17 NET171 NET170 WL BIT_B_17 SRAM_CELL_G1 
XI17 BIT_16 NET176 NET175 WL BIT_B_16 SRAM_CELL_G1 
XI16 BIT_15 NET181 NET180 WL BIT_B_15 SRAM_CELL_G1 
XI15 BIT_14 NET186 NET185 WL BIT_B_14 SRAM_CELL_G1 
XI14 BIT_13 NET191 NET190 WL BIT_B_13 SRAM_CELL_G1 
XI13 BIT_12 NET196 NET195 WL BIT_B_12 SRAM_CELL_G1 
XI12 BIT_11 NET201 NET200 WL BIT_B_11 SRAM_CELL_G1 
XI11 BIT_10 NET206 NET205 WL BIT_B_10 SRAM_CELL_G1 
XI10 BIT_9 NET211 NET210 WL BIT_B_9 SRAM_CELL_G1 
XI9 BIT_8 NET216 NET215 WL BIT_B_8 SRAM_CELL_G1 
XI8 BIT_7 NET221 NET220 WL BIT_B_7 SRAM_CELL_G1 
XI7 BIT_6 NET226 NET225 WL BIT_B_6 SRAM_CELL_G1 
XI6 BIT_5 NET231 NET230 WL BIT_B_5 SRAM_CELL_G1 
XI5 BIT_4 NET236 NET235 WL BIT_B_4 SRAM_CELL_G1 
XI4 BIT_3 NET241 NET240 WL BIT_B_3 SRAM_CELL_G1 
XI3 BIT_2 NET246 NET245 WL BIT_B_2 SRAM_CELL_G1 
XI2 BIT_1 NET251 NET250 WL BIT_B_1 SRAM_CELL_G1 
XI1 BIT_0 NET256 NET255 WL BIT_B_0 SRAM_CELL_G1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SRAM_CELL32_G3 
* FILE NAME: SRAM2_REG10_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: REG10.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:36 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   IN<0> = IN_0
*                   IN<1> = IN_1
*                   IN<2> = IN_2
*                   IN<3> = IN_3
*                   IN<4> = IN_4
*                   IN<5> = IN_5
*                   IN<6> = IN_6
*                   IN<7> = IN_7
*                   IN<8> = IN_8
*                   IN<9> = IN_9
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
*                   OUT<3> = OUT_3
*                   OUT<4> = OUT_4
*                   OUT<5> = OUT_5
*                   OUT<6> = OUT_6
*                   OUT<7> = OUT_7
*                   OUT<8> = OUT_8
*                   OUT<9> = OUT_9
.SUBCKT REG10_G21 CLK IN_0 IN_1 IN_2 IN_3 IN_4 IN_5 IN_6 IN_7 IN_8 IN_9 OUT_0 
+OUT_1 OUT_2 OUT_3 OUT_4 OUT_5 OUT_6 OUT_7 OUT_8 OUT_9 
XI9 CLK IN_9 OUT_9 DFFPOSX1_G6 
XI8 CLK IN_8 OUT_8 DFFPOSX1_G6 
XI7 CLK IN_7 OUT_7 DFFPOSX1_G6 
XI6 CLK IN_6 OUT_6 DFFPOSX1_G6 
XI5 CLK IN_5 OUT_5 DFFPOSX1_G6 
XI4 CLK IN_4 OUT_4 DFFPOSX1_G6 
XI3 CLK IN_3 OUT_3 DFFPOSX1_G6 
XI2 CLK IN_2 OUT_2 DFFPOSX1_G6 
XI1 CLK IN_1 OUT_1 DFFPOSX1_G6 
XI0 CLK IN_0 OUT_0 DFFPOSX1_G6 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS REG10_G21 
* FILE NAME: SRAM2_SAMP_CELL32_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SAMP_CELL32.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:43 2007.
   
* TERMINAL MAPPING: BIT<0> = BIT_0
*                   BIT<1> = BIT_1
*                   BIT<2> = BIT_2
*                   BIT<3> = BIT_3
*                   BIT<4> = BIT_4
*                   BIT<5> = BIT_5
*                   BIT<6> = BIT_6
*                   BIT<7> = BIT_7
*                   BIT<8> = BIT_8
*                   BIT<9> = BIT_9
*                   BIT<10> = BIT_10
*                   BIT<11> = BIT_11
*                   BIT<12> = BIT_12
*                   BIT<13> = BIT_13
*                   BIT<14> = BIT_14
*                   BIT<15> = BIT_15
*                   BIT<16> = BIT_16
*                   BIT<17> = BIT_17
*                   BIT<18> = BIT_18
*                   BIT<19> = BIT_19
*                   BIT<20> = BIT_20
*                   BIT<21> = BIT_21
*                   BIT<22> = BIT_22
*                   BIT<23> = BIT_23
*                   BIT<24> = BIT_24
*                   BIT<25> = BIT_25
*                   BIT<26> = BIT_26
*                   BIT<27> = BIT_27
*                   BIT<28> = BIT_28
*                   BIT<29> = BIT_29
*                   BIT<30> = BIT_30
*                   BIT<31> = BIT_31
*                   BIT_B<0> = BIT_B_0
*                   BIT_B<1> = BIT_B_1
*                   BIT_B<2> = BIT_B_2
*                   BIT_B<3> = BIT_B_3
*                   BIT_B<4> = BIT_B_4
*                   BIT_B<5> = BIT_B_5
*                   BIT_B<6> = BIT_B_6
*                   BIT_B<7> = BIT_B_7
*                   BIT_B<8> = BIT_B_8
*                   BIT_B<9> = BIT_B_9
*                   BIT_B<10> = BIT_B_10
*                   BIT_B<11> = BIT_B_11
*                   BIT_B<12> = BIT_B_12
*                   BIT_B<13> = BIT_B_13
*                   BIT_B<14> = BIT_B_14
*                   BIT_B<15> = BIT_B_15
*                   BIT_B<16> = BIT_B_16
*                   BIT_B<17> = BIT_B_17
*                   BIT_B<18> = BIT_B_18
*                   BIT_B<19> = BIT_B_19
*                   BIT_B<20> = BIT_B_20
*                   BIT_B<21> = BIT_B_21
*                   BIT_B<22> = BIT_B_22
*                   BIT_B<23> = BIT_B_23
*                   BIT_B<24> = BIT_B_24
*                   BIT_B<25> = BIT_B_25
*                   BIT_B<26> = BIT_B_26
*                   BIT_B<27> = BIT_B_27
*                   BIT_B<28> = BIT_B_28
*                   BIT_B<29> = BIT_B_29
*                   BIT_B<30> = BIT_B_30
*                   BIT_B<31> = BIT_B_31
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
*                   OUT<3> = OUT_3
*                   OUT<4> = OUT_4
*                   OUT<5> = OUT_5
*                   OUT<6> = OUT_6
*                   OUT<7> = OUT_7
*                   OUT<8> = OUT_8
*                   OUT<9> = OUT_9
*                   OUT<10> = OUT_10
*                   OUT<11> = OUT_11
*                   OUT<12> = OUT_12
*                   OUT<13> = OUT_13
*                   OUT<14> = OUT_14
*                   OUT<15> = OUT_15
*                   OUT<16> = OUT_16
*                   OUT<17> = OUT_17
*                   OUT<18> = OUT_18
*                   OUT<19> = OUT_19
*                   OUT<20> = OUT_20
*                   OUT<21> = OUT_21
*                   OUT<22> = OUT_22
*                   OUT<23> = OUT_23
*                   OUT<24> = OUT_24
*                   OUT<25> = OUT_25
*                   OUT<26> = OUT_26
*                   OUT<27> = OUT_27
*                   OUT<28> = OUT_28
*                   OUT<29> = OUT_29
*                   OUT<30> = OUT_30
*                   OUT<31> = OUT_31
*                   OUT_B<0> = OUT_B_0
*                   OUT_B<1> = OUT_B_1
*                   OUT_B<2> = OUT_B_2
*                   OUT_B<3> = OUT_B_3
*                   OUT_B<4> = OUT_B_4
*                   OUT_B<5> = OUT_B_5
*                   OUT_B<6> = OUT_B_6
*                   OUT_B<7> = OUT_B_7
*                   OUT_B<8> = OUT_B_8
*                   OUT_B<9> = OUT_B_9
*                   OUT_B<10> = OUT_B_10
*                   OUT_B<11> = OUT_B_11
*                   OUT_B<12> = OUT_B_12
*                   OUT_B<13> = OUT_B_13
*                   OUT_B<14> = OUT_B_14
*                   OUT_B<15> = OUT_B_15
*                   OUT_B<16> = OUT_B_16
*                   OUT_B<17> = OUT_B_17
*                   OUT_B<18> = OUT_B_18
*                   OUT_B<19> = OUT_B_19
*                   OUT_B<20> = OUT_B_20
*                   OUT_B<21> = OUT_B_21
*                   OUT_B<22> = OUT_B_22
*                   OUT_B<23> = OUT_B_23
*                   OUT_B<24> = OUT_B_24
*                   OUT_B<25> = OUT_B_25
*                   OUT_B<26> = OUT_B_26
*                   OUT_B<27> = OUT_B_27
*                   OUT_B<28> = OUT_B_28
*                   OUT_B<29> = OUT_B_29
*                   OUT_B<30> = OUT_B_30
*                   OUT_B<31> = OUT_B_31
*                   READ_EN = READ_EN
.SUBCKT SAMP_CELL32_G26 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 BIT_8 
+BIT_9 BIT_10 BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 BIT_19 
+BIT_20 BIT_21 BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 BIT_30 
+BIT_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 
+BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 
+BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 
+BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 BIT_B_29 BIT_B_30 BIT_B_31 OUT_0 OUT_1 
+OUT_2 OUT_3 OUT_4 OUT_5 OUT_6 OUT_7 OUT_8 OUT_9 OUT_10 OUT_11 OUT_12 OUT_13 
+OUT_14 OUT_15 OUT_16 OUT_17 OUT_18 OUT_19 OUT_20 OUT_21 OUT_22 OUT_23 OUT_24 
+OUT_25 OUT_26 OUT_27 OUT_28 OUT_29 OUT_30 OUT_31 OUT_B_0 OUT_B_1 OUT_B_2 
+OUT_B_3 OUT_B_4 OUT_B_5 OUT_B_6 OUT_B_7 OUT_B_8 OUT_B_9 OUT_B_10 OUT_B_11 
+OUT_B_12 OUT_B_13 OUT_B_14 OUT_B_15 OUT_B_16 OUT_B_17 OUT_B_18 OUT_B_19 
+OUT_B_20 OUT_B_21 OUT_B_22 OUT_B_23 OUT_B_24 OUT_B_25 OUT_B_26 OUT_B_27 
+OUT_B_28 OUT_B_29 OUT_B_30 OUT_B_31 READ_EN 
XI1 BIT_1 OUT_1 BIT_B_1 OUT_B_1 READ_EN SAMP_CELL_G12 
XI0 BIT_0 OUT_0 BIT_B_0 OUT_B_0 READ_EN SAMP_CELL_G12 
XI31 BIT_31 OUT_31 BIT_B_31 OUT_B_31 READ_EN SAMP_CELL_G12 
XI30 BIT_30 OUT_30 BIT_B_30 OUT_B_30 READ_EN SAMP_CELL_G12 
XI29 BIT_29 OUT_29 BIT_B_29 OUT_B_29 READ_EN SAMP_CELL_G12 
XI28 BIT_28 OUT_28 BIT_B_28 OUT_B_28 READ_EN SAMP_CELL_G12 
XI27 BIT_27 OUT_27 BIT_B_27 OUT_B_27 READ_EN SAMP_CELL_G12 
XI26 BIT_26 OUT_26 BIT_B_26 OUT_B_26 READ_EN SAMP_CELL_G12 
XI25 BIT_25 OUT_25 BIT_B_25 OUT_B_25 READ_EN SAMP_CELL_G12 
XI24 BIT_24 OUT_24 BIT_B_24 OUT_B_24 READ_EN SAMP_CELL_G12 
XI23 BIT_23 OUT_23 BIT_B_23 OUT_B_23 READ_EN SAMP_CELL_G12 
XI22 BIT_22 OUT_22 BIT_B_22 OUT_B_22 READ_EN SAMP_CELL_G12 
XI21 BIT_21 OUT_21 BIT_B_21 OUT_B_21 READ_EN SAMP_CELL_G12 
XI20 BIT_20 OUT_20 BIT_B_20 OUT_B_20 READ_EN SAMP_CELL_G12 
XI19 BIT_19 OUT_19 BIT_B_19 OUT_B_19 READ_EN SAMP_CELL_G12 
XI18 BIT_18 OUT_18 BIT_B_18 OUT_B_18 READ_EN SAMP_CELL_G12 
XI17 BIT_17 OUT_17 BIT_B_17 OUT_B_17 READ_EN SAMP_CELL_G12 
XI16 BIT_16 OUT_16 BIT_B_16 OUT_B_16 READ_EN SAMP_CELL_G12 
XI15 BIT_15 OUT_15 BIT_B_15 OUT_B_15 READ_EN SAMP_CELL_G12 
XI14 BIT_14 OUT_14 BIT_B_14 OUT_B_14 READ_EN SAMP_CELL_G12 
XI13 BIT_13 OUT_13 BIT_B_13 OUT_B_13 READ_EN SAMP_CELL_G12 
XI12 BIT_12 OUT_12 BIT_B_12 OUT_B_12 READ_EN SAMP_CELL_G12 
XI11 BIT_11 OUT_11 BIT_B_11 OUT_B_11 READ_EN SAMP_CELL_G12 
XI10 BIT_10 OUT_10 BIT_B_10 OUT_B_10 READ_EN SAMP_CELL_G12 
XI9 BIT_9 OUT_9 BIT_B_9 OUT_B_9 READ_EN SAMP_CELL_G12 
XI8 BIT_8 OUT_8 BIT_B_8 OUT_B_8 READ_EN SAMP_CELL_G12 
XI7 BIT_7 OUT_7 BIT_B_7 OUT_B_7 READ_EN SAMP_CELL_G12 
XI6 BIT_6 OUT_6 BIT_B_6 OUT_B_6 READ_EN SAMP_CELL_G12 
XI5 BIT_5 OUT_5 BIT_B_5 OUT_B_5 READ_EN SAMP_CELL_G12 
XI4 BIT_4 OUT_4 BIT_B_4 OUT_B_4 READ_EN SAMP_CELL_G12 
XI3 BIT_3 OUT_3 BIT_B_3 OUT_B_3 READ_EN SAMP_CELL_G12 
XI2 BIT_2 OUT_2 BIT_B_2 OUT_B_2 READ_EN SAMP_CELL_G12 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SAMP_CELL32_G26 
* FILE NAME: SRAM2_WRITE_CELL32_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: WRITE_CELL32.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:43 2007.
   
* TERMINAL MAPPING: BT1<0> = BT1_0
*                   BT1<1> = BT1_1
*                   BT1<2> = BT1_2
*                   BT1<3> = BT1_3
*                   BT1<4> = BT1_4
*                   BT1<5> = BT1_5
*                   BT1<6> = BT1_6
*                   BT1<7> = BT1_7
*                   BT1<8> = BT1_8
*                   BT1<9> = BT1_9
*                   BT1<10> = BT1_10
*                   BT1<11> = BT1_11
*                   BT1<12> = BT1_12
*                   BT1<13> = BT1_13
*                   BT1<14> = BT1_14
*                   BT1<15> = BT1_15
*                   BT1<16> = BT1_16
*                   BT1<17> = BT1_17
*                   BT1<18> = BT1_18
*                   BT1<19> = BT1_19
*                   BT1<20> = BT1_20
*                   BT1<21> = BT1_21
*                   BT1<22> = BT1_22
*                   BT1<23> = BT1_23
*                   BT1<24> = BT1_24
*                   BT1<25> = BT1_25
*                   BT1<26> = BT1_26
*                   BT1<27> = BT1_27
*                   BT1<28> = BT1_28
*                   BT1<29> = BT1_29
*                   BT1<30> = BT1_30
*                   BT1<31> = BT1_31
*                   BT2<0> = BT2_0
*                   BT2<1> = BT2_1
*                   BT2<2> = BT2_2
*                   BT2<3> = BT2_3
*                   BT2<4> = BT2_4
*                   BT2<5> = BT2_5
*                   BT2<6> = BT2_6
*                   BT2<7> = BT2_7
*                   BT2<8> = BT2_8
*                   BT2<9> = BT2_9
*                   BT2<10> = BT2_10
*                   BT2<11> = BT2_11
*                   BT2<12> = BT2_12
*                   BT2<13> = BT2_13
*                   BT2<14> = BT2_14
*                   BT2<15> = BT2_15
*                   BT2<16> = BT2_16
*                   BT2<17> = BT2_17
*                   BT2<18> = BT2_18
*                   BT2<19> = BT2_19
*                   BT2<20> = BT2_20
*                   BT2<21> = BT2_21
*                   BT2<22> = BT2_22
*                   BT2<23> = BT2_23
*                   BT2<24> = BT2_24
*                   BT2<25> = BT2_25
*                   BT2<26> = BT2_26
*                   BT2<27> = BT2_27
*                   BT2<28> = BT2_28
*                   BT2<29> = BT2_29
*                   BT2<30> = BT2_30
*                   BT2<31> = BT2_31
*                   BTB1<0> = BTB1_0
*                   BTB1<1> = BTB1_1
*                   BTB1<2> = BTB1_2
*                   BTB1<3> = BTB1_3
*                   BTB1<4> = BTB1_4
*                   BTB1<5> = BTB1_5
*                   BTB1<6> = BTB1_6
*                   BTB1<7> = BTB1_7
*                   BTB1<8> = BTB1_8
*                   BTB1<9> = BTB1_9
*                   BTB1<10> = BTB1_10
*                   BTB1<11> = BTB1_11
*                   BTB1<12> = BTB1_12
*                   BTB1<13> = BTB1_13
*                   BTB1<14> = BTB1_14
*                   BTB1<15> = BTB1_15
*                   BTB1<16> = BTB1_16
*                   BTB1<17> = BTB1_17
*                   BTB1<18> = BTB1_18
*                   BTB1<19> = BTB1_19
*                   BTB1<20> = BTB1_20
*                   BTB1<21> = BTB1_21
*                   BTB1<22> = BTB1_22
*                   BTB1<23> = BTB1_23
*                   BTB1<24> = BTB1_24
*                   BTB1<25> = BTB1_25
*                   BTB1<26> = BTB1_26
*                   BTB1<27> = BTB1_27
*                   BTB1<28> = BTB1_28
*                   BTB1<29> = BTB1_29
*                   BTB1<30> = BTB1_30
*                   BTB1<31> = BTB1_31
*                   BTB2<0> = BTB2_0
*                   BTB2<1> = BTB2_1
*                   BTB2<2> = BTB2_2
*                   BTB2<3> = BTB2_3
*                   BTB2<4> = BTB2_4
*                   BTB2<5> = BTB2_5
*                   BTB2<6> = BTB2_6
*                   BTB2<7> = BTB2_7
*                   BTB2<8> = BTB2_8
*                   BTB2<9> = BTB2_9
*                   BTB2<10> = BTB2_10
*                   BTB2<11> = BTB2_11
*                   BTB2<12> = BTB2_12
*                   BTB2<13> = BTB2_13
*                   BTB2<14> = BTB2_14
*                   BTB2<15> = BTB2_15
*                   BTB2<16> = BTB2_16
*                   BTB2<17> = BTB2_17
*                   BTB2<18> = BTB2_18
*                   BTB2<19> = BTB2_19
*                   BTB2<20> = BTB2_20
*                   BTB2<21> = BTB2_21
*                   BTB2<22> = BTB2_22
*                   BTB2<23> = BTB2_23
*                   BTB2<24> = BTB2_24
*                   BTB2<25> = BTB2_25
*                   BTB2<26> = BTB2_26
*                   BTB2<27> = BTB2_27
*                   BTB2<28> = BTB2_28
*                   BTB2<29> = BTB2_29
*                   BTB2<30> = BTB2_30
*                   BTB2<31> = BTB2_31
*                   DATA<0> = DATA_0
*                   DATA<1> = DATA_1
*                   DATA<2> = DATA_2
*                   DATA<3> = DATA_3
*                   DATA<4> = DATA_4
*                   DATA<5> = DATA_5
*                   DATA<6> = DATA_6
*                   DATA<7> = DATA_7
*                   DATA<8> = DATA_8
*                   DATA<9> = DATA_9
*                   DATA<10> = DATA_10
*                   DATA<11> = DATA_11
*                   DATA<12> = DATA_12
*                   DATA<13> = DATA_13
*                   DATA<14> = DATA_14
*                   DATA<15> = DATA_15
*                   DATA<16> = DATA_16
*                   DATA<17> = DATA_17
*                   DATA<18> = DATA_18
*                   DATA<19> = DATA_19
*                   DATA<20> = DATA_20
*                   DATA<21> = DATA_21
*                   DATA<22> = DATA_22
*                   DATA<23> = DATA_23
*                   DATA<24> = DATA_24
*                   DATA<25> = DATA_25
*                   DATA<26> = DATA_26
*                   DATA<27> = DATA_27
*                   DATA<28> = DATA_28
*                   DATA<29> = DATA_29
*                   DATA<30> = DATA_30
*                   DATA<31> = DATA_31
*                   DATA_B<0> = DATA_B_0
*                   DATA_B<1> = DATA_B_1
*                   DATA_B<2> = DATA_B_2
*                   DATA_B<3> = DATA_B_3
*                   DATA_B<4> = DATA_B_4
*                   DATA_B<5> = DATA_B_5
*                   DATA_B<6> = DATA_B_6
*                   DATA_B<7> = DATA_B_7
*                   DATA_B<8> = DATA_B_8
*                   DATA_B<9> = DATA_B_9
*                   DATA_B<10> = DATA_B_10
*                   DATA_B<11> = DATA_B_11
*                   DATA_B<12> = DATA_B_12
*                   DATA_B<13> = DATA_B_13
*                   DATA_B<14> = DATA_B_14
*                   DATA_B<15> = DATA_B_15
*                   DATA_B<16> = DATA_B_16
*                   DATA_B<17> = DATA_B_17
*                   DATA_B<18> = DATA_B_18
*                   DATA_B<19> = DATA_B_19
*                   DATA_B<20> = DATA_B_20
*                   DATA_B<21> = DATA_B_21
*                   DATA_B<22> = DATA_B_22
*                   DATA_B<23> = DATA_B_23
*                   DATA_B<24> = DATA_B_24
*                   DATA_B<25> = DATA_B_25
*                   DATA_B<26> = DATA_B_26
*                   DATA_B<27> = DATA_B_27
*                   DATA_B<28> = DATA_B_28
*                   DATA_B<29> = DATA_B_29
*                   DATA_B<30> = DATA_B_30
*                   DATA_B<31> = DATA_B_31
*                   PRE = PRE
*                   WRITE_EN = WRITE_EN
.SUBCKT WRITE_CELL32_G25 BT1_0 BT1_1 BT1_2 BT1_3 BT1_4 BT1_5 BT1_6 BT1_7 BT1_8 
+BT1_9 BT1_10 BT1_11 BT1_12 BT1_13 BT1_14 BT1_15 BT1_16 BT1_17 BT1_18 BT1_19 
+BT1_20 BT1_21 BT1_22 BT1_23 BT1_24 BT1_25 BT1_26 BT1_27 BT1_28 BT1_29 BT1_30 
+BT1_31 BT2_0 BT2_1 BT2_2 BT2_3 BT2_4 BT2_5 BT2_6 BT2_7 BT2_8 BT2_9 BT2_10 
+BT2_11 BT2_12 BT2_13 BT2_14 BT2_15 BT2_16 BT2_17 BT2_18 BT2_19 BT2_20 BT2_21 
+BT2_22 BT2_23 BT2_24 BT2_25 BT2_26 BT2_27 BT2_28 BT2_29 BT2_30 BT2_31 BTB1_0 
+BTB1_1 BTB1_2 BTB1_3 BTB1_4 BTB1_5 BTB1_6 BTB1_7 BTB1_8 BTB1_9 BTB1_10 BTB1_11 
+BTB1_12 BTB1_13 BTB1_14 BTB1_15 BTB1_16 BTB1_17 BTB1_18 BTB1_19 BTB1_20 
+BTB1_21 BTB1_22 BTB1_23 BTB1_24 BTB1_25 BTB1_26 BTB1_27 BTB1_28 BTB1_29 
+BTB1_30 BTB1_31 BTB2_0 BTB2_1 BTB2_2 BTB2_3 BTB2_4 BTB2_5 BTB2_6 BTB2_7 BTB2_8 
+BTB2_9 BTB2_10 BTB2_11 BTB2_12 BTB2_13 BTB2_14 BTB2_15 BTB2_16 BTB2_17 BTB2_18 
+BTB2_19 BTB2_20 BTB2_21 BTB2_22 BTB2_23 BTB2_24 BTB2_25 BTB2_26 BTB2_27 
+BTB2_28 BTB2_29 BTB2_30 BTB2_31 DATA_0 DATA_1 DATA_2 DATA_3 DATA_4 DATA_5 
+DATA_6 DATA_7 DATA_8 DATA_9 DATA_10 DATA_11 DATA_12 DATA_13 DATA_14 DATA_15 
+DATA_16 DATA_17 DATA_18 DATA_19 DATA_20 DATA_21 DATA_22 DATA_23 DATA_24 
+DATA_25 DATA_26 DATA_27 DATA_28 DATA_29 DATA_30 DATA_31 DATA_B_0 DATA_B_1 
+DATA_B_2 DATA_B_3 DATA_B_4 DATA_B_5 DATA_B_6 DATA_B_7 DATA_B_8 DATA_B_9 
+DATA_B_10 DATA_B_11 DATA_B_12 DATA_B_13 DATA_B_14 DATA_B_15 DATA_B_16 
+DATA_B_17 DATA_B_18 DATA_B_19 DATA_B_20 DATA_B_21 DATA_B_22 DATA_B_23 
+DATA_B_24 DATA_B_25 DATA_B_26 DATA_B_27 DATA_B_28 DATA_B_29 DATA_B_30 
+DATA_B_31 PRE WRITE_EN 
XI31 BT1_31 BT2_31 BTB1_31 BTB2_31 DATA_31 PRE DATA_B_31 WRITE_EN 
+WRITE_CELL_G11 
XI30 BT1_30 BT2_30 BTB1_30 BTB2_30 DATA_30 PRE DATA_B_30 WRITE_EN 
+WRITE_CELL_G11 
XI29 BT1_29 BT2_29 BTB1_29 BTB2_29 DATA_29 PRE DATA_B_29 WRITE_EN 
+WRITE_CELL_G11 
XI28 BT1_28 BT2_28 BTB1_28 BTB2_28 DATA_28 PRE DATA_B_28 WRITE_EN 
+WRITE_CELL_G11 
XI27 BT1_27 BT2_27 BTB1_27 BTB2_27 DATA_27 PRE DATA_B_27 WRITE_EN 
+WRITE_CELL_G11 
XI26 BT1_26 BT2_26 BTB1_26 BTB2_26 DATA_26 PRE DATA_B_26 WRITE_EN 
+WRITE_CELL_G11 
XI25 BT1_25 BT2_25 BTB1_25 BTB2_25 DATA_25 PRE DATA_B_25 WRITE_EN 
+WRITE_CELL_G11 
XI24 BT1_24 BT2_24 BTB1_24 BTB2_24 DATA_24 PRE DATA_B_24 WRITE_EN 
+WRITE_CELL_G11 
XI23 BT1_23 BT2_23 BTB1_23 BTB2_23 DATA_23 PRE DATA_B_23 WRITE_EN 
+WRITE_CELL_G11 
XI22 BT1_22 BT2_22 BTB1_22 BTB2_22 DATA_22 PRE DATA_B_22 WRITE_EN 
+WRITE_CELL_G11 
XI21 BT1_21 BT2_21 BTB1_21 BTB2_21 DATA_21 PRE DATA_B_21 WRITE_EN 
+WRITE_CELL_G11 
XI20 BT1_20 BT2_20 BTB1_20 BTB2_20 DATA_20 PRE DATA_B_20 WRITE_EN 
+WRITE_CELL_G11 
XI19 BT1_19 BT2_19 BTB1_19 BTB2_19 DATA_19 PRE DATA_B_19 WRITE_EN 
+WRITE_CELL_G11 
XI18 BT1_18 BT2_18 BTB1_18 BTB2_18 DATA_18 PRE DATA_B_18 WRITE_EN 
+WRITE_CELL_G11 
XI17 BT1_17 BT2_17 BTB1_17 BTB2_17 DATA_17 PRE DATA_B_17 WRITE_EN 
+WRITE_CELL_G11 
XI16 BT1_16 BT2_16 BTB1_16 BTB2_16 DATA_16 PRE DATA_B_16 WRITE_EN 
+WRITE_CELL_G11 
XI15 BT1_15 BT2_15 BTB1_15 BTB2_15 DATA_15 PRE DATA_B_15 WRITE_EN 
+WRITE_CELL_G11 
XI14 BT1_14 BT2_14 BTB1_14 BTB2_14 DATA_14 PRE DATA_B_14 WRITE_EN 
+WRITE_CELL_G11 
XI13 BT1_13 BT2_13 BTB1_13 BTB2_13 DATA_13 PRE DATA_B_13 WRITE_EN 
+WRITE_CELL_G11 
XI12 BT1_12 BT2_12 BTB1_12 BTB2_12 DATA_12 PRE DATA_B_12 WRITE_EN 
+WRITE_CELL_G11 
XI11 BT1_11 BT2_11 BTB1_11 BTB2_11 DATA_11 PRE DATA_B_11 WRITE_EN 
+WRITE_CELL_G11 
XI10 BT1_10 BT2_10 BTB1_10 BTB2_10 DATA_10 PRE DATA_B_10 WRITE_EN 
+WRITE_CELL_G11 
XI9 BT1_9 BT2_9 BTB1_9 BTB2_9 DATA_9 PRE DATA_B_9 WRITE_EN WRITE_CELL_G11 
XI8 BT1_8 BT2_8 BTB1_8 BTB2_8 DATA_8 PRE DATA_B_8 WRITE_EN WRITE_CELL_G11 
XI7 BT1_7 BT2_7 BTB1_7 BTB2_7 DATA_7 PRE DATA_B_7 WRITE_EN WRITE_CELL_G11 
XI6 BT1_6 BT2_6 BTB1_6 BTB2_6 DATA_6 PRE DATA_B_6 WRITE_EN WRITE_CELL_G11 
XI5 BT1_5 BT2_5 BTB1_5 BTB2_5 DATA_5 PRE DATA_B_5 WRITE_EN WRITE_CELL_G11 
XI4 BT1_4 BT2_4 BTB1_4 BTB2_4 DATA_4 PRE DATA_B_4 WRITE_EN WRITE_CELL_G11 
XI3 BT1_3 BT2_3 BTB1_3 BTB2_3 DATA_3 PRE DATA_B_3 WRITE_EN WRITE_CELL_G11 
XI2 BT1_2 BT2_2 BTB1_2 BTB2_2 DATA_2 PRE DATA_B_2 WRITE_EN WRITE_CELL_G11 
XI1 BT1_1 BT2_1 BTB1_1 BTB2_1 DATA_1 PRE DATA_B_1 WRITE_EN WRITE_CELL_G11 
XI0 BT1_0 BT2_0 BTB1_0 BTB2_0 DATA_0 PRE DATA_B_0 WRITE_EN WRITE_CELL_G11 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS WRITE_CELL32_G25 
* FILE NAME: SRAM2_WRITE_CELL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: WRITE_CELL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:43 2007.
   
* TERMINAL MAPPING: BT1 = BT1
*                   BT2 = BT2
*                   BTB1 = BTB1
*                   BTB2 = BTB2
*                   DATA = DATA
*                   PRE = PRE
*                   DATA_BAR = DATA_BAR
*                   WRITE_EN = WRITE_EN
.SUBCKT WRITE_CELL_G11 BT1 BT2 BTB1 BTB2 DATA PRE DATA_BAR WRITE_EN 
M5 BTB1 PRE VDD! VDD!  PFET  L=200E-9 W=12E-6 AD=+6.00000000E-12 
+AS=+6.00000000E-12 PD=+2.50000000E-05 PS=+2.50000000E-05 NRD=+4.16666667E-02 
+NRS=+4.16666667E-02 M=1.0 
M1 BT1 PRE VDD! VDD!  PFET  L=200E-9 W=12E-6 AD=+6.00000000E-12 
+AS=+6.00000000E-12 PD=+2.50000000E-05 PS=+2.50000000E-05 NRD=+4.16666667E-02 
+NRS=+4.16666667E-02 M=1.0 
M4 NET17 DATA 0 0  NFET  L=200E-9 W=3.4E-6 AD=+1.70000000E-12 
+AS=+1.70000000E-12 PD=+7.80000000E-06 PS=+7.80000000E-06 NRD=+1.47058824E-01 
+NRS=+1.47058824E-01 M=1.0 
M3 BTB2 WRITE_EN NET17 0  NFET  L=200E-9 W=3.4E-6 AD=+1.70000000E-12 
+AS=+1.70000000E-12 PD=+7.80000000E-06 PS=+7.80000000E-06 NRD=+1.47058824E-01 
+NRS=+1.47058824E-01 M=1.0 
M2 BT2 WRITE_EN NET26 0  NFET  L=200E-9 W=3.4E-6 AD=+1.70000000E-12 
+AS=+1.70000000E-12 PD=+7.80000000E-06 PS=+7.80000000E-06 NRD=+1.47058824E-01 
+NRS=+1.47058824E-01 M=1.0 
M0 NET26 DATA_BAR 0 0  NFET  L=200E-9 W=3.4E-6 AD=+1.70000000E-12 
+AS=+1.70000000E-12 PD=+7.80000000E-06 PS=+7.80000000E-06 NRD=+1.47058824E-01 
+NRS=+1.47058824E-01 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS WRITE_CELL_G11 
* FILE NAME: SRAM2_RDEC3TO8A_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: RDEC3TO8A.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:35 2007.
   
* TERMINAL MAPPING: RDECO<0> = RDECO_0
*                   RDECO<1> = RDECO_1
*                   RDECO<2> = RDECO_2
*                   RDECO<3> = RDECO_3
*                   RDECO<4> = RDECO_4
*                   RDECO<5> = RDECO_5
*                   RDECO<6> = RDECO_6
*                   RDECO<7> = RDECO_7
*                   RI<0> = RI_0
*                   RI<1> = RI_1
*                   RI<2> = RI_2
*                   RIB<0> = RIB_0
*                   RIB<1> = RIB_1
*                   RIB<2> = RIB_2
*                   TOP = TOP
.SUBCKT RDEC3TO8A_G4 RDECO_0 RDECO_1 RDECO_2 RDECO_3 RDECO_4 RDECO_5 RDECO_6 
+RDECO_7 RI_0 RI_1 RI_2 RIB_0 RIB_1 RIB_2 TOP 
M37 NET0174 RIB_2 TOP VDD!  PFET  L=200E-9 W=9.6E-6 AD=+4.80000000E-12 
+AS=+4.80000000E-12 PD=+2.02000000E-05 PS=+2.02000000E-05 NRD=+5.20833333E-02 
+NRS=+5.20833333E-02 M=1.0 
M36 NET0175 RI_2 TOP VDD!  PFET  L=200E-9 W=9.6E-6 AD=+4.80000000E-12 
+AS=+4.80000000E-12 PD=+2.02000000E-05 PS=+2.02000000E-05 NRD=+5.20833333E-02 
+NRS=+5.20833333E-02 M=1.0 
M28 RDECO_1 RIB_0 NET056 VDD!  PFET  L=200E-9 W=2.4E-6 AD=+1.20000000E-12 
+AS=+1.20000000E-12 PD=+5.80000000E-06 PS=+5.80000000E-06 NRD=+2.08333333E-01 
+NRS=+2.08333333E-01 M=1.0 
M29 RDECO_3 RIB_0 NET068 VDD!  PFET  L=200E-9 W=2.4E-6 AD=+1.20000000E-12 
+AS=+1.20000000E-12 PD=+5.80000000E-06 PS=+5.80000000E-06 NRD=+2.08333333E-01 
+NRS=+2.08333333E-01 M=1.0 
M30 RDECO_5 RIB_0 NET050 VDD!  PFET  L=200E-9 W=2.4E-6 AD=+1.20000000E-12 
+AS=+1.20000000E-12 PD=+5.80000000E-06 PS=+5.80000000E-06 NRD=+2.08333333E-01 
+NRS=+2.08333333E-01 M=1.0 
M31 RDECO_7 RIB_0 NET062 VDD!  PFET  L=200E-9 W=2.4E-6 AD=+1.20000000E-12 
+AS=+1.20000000E-12 PD=+5.80000000E-06 PS=+5.80000000E-06 NRD=+2.08333333E-01 
+NRS=+2.08333333E-01 M=1.0 
M8 RDECO_0 RI_0 NET056 VDD!  PFET  L=200E-9 W=2.4E-6 AD=+1.20000000E-12 
+AS=+1.20000000E-12 PD=+5.80000000E-06 PS=+5.80000000E-06 NRD=+2.08333333E-01 
+NRS=+2.08333333E-01 M=1.0 
M27 RDECO_6 RI_0 NET062 VDD!  PFET  L=200E-9 W=2.4E-6 AD=+1.20000000E-12 
+AS=+1.20000000E-12 PD=+5.80000000E-06 PS=+5.80000000E-06 NRD=+2.08333333E-01 
+NRS=+2.08333333E-01 M=1.0 
M32 NET056 RI_1 NET0175 VDD!  PFET  L=200E-9 W=4.8E-6 AD=+2.40000000E-12 
+AS=+2.40000000E-12 PD=+1.06000000E-05 PS=+1.06000000E-05 NRD=+1.04166667E-01 
+NRS=+1.04166667E-01 M=1.0 
M33 NET050 RI_1 NET0174 VDD!  PFET  L=200E-9 W=4.8E-6 AD=+2.40000000E-12 
+AS=+2.40000000E-12 PD=+1.06000000E-05 PS=+1.06000000E-05 NRD=+1.04166667E-01 
+NRS=+1.04166667E-01 M=1.0 
M34 NET068 RIB_1 NET0175 VDD!  PFET  L=200E-9 W=4.8E-6 AD=+2.40000000E-12 
+AS=+2.40000000E-12 PD=+1.06000000E-05 PS=+1.06000000E-05 NRD=+1.04166667E-01 
+NRS=+1.04166667E-01 M=1.0 
M35 NET062 RIB_1 NET0174 VDD!  PFET  L=200E-9 W=4.8E-6 AD=+2.40000000E-12 
+AS=+2.40000000E-12 PD=+1.06000000E-05 PS=+1.06000000E-05 NRD=+1.04166667E-01 
+NRS=+1.04166667E-01 M=1.0 
M26 RDECO_4 RI_0 NET050 VDD!  PFET  L=200E-9 W=2.4E-6 AD=+1.20000000E-12 
+AS=+1.20000000E-12 PD=+5.80000000E-06 PS=+5.80000000E-06 NRD=+2.08333333E-01 
+NRS=+2.08333333E-01 M=1.0 
M25 RDECO_2 RI_0 NET068 VDD!  PFET  L=200E-9 W=2.4E-6 AD=+1.20000000E-12 
+AS=+1.20000000E-12 PD=+5.80000000E-06 PS=+5.80000000E-06 NRD=+2.08333333E-01 
+NRS=+2.08333333E-01 M=1.0 
M24 RDECO_0 RI_1 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M23 RDECO_7 RIB_2 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M22 RDECO_6 RIB_2 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M21 RDECO_5 RIB_2 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M20 RDECO_4 RIB_2 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M19 RDECO_3 RI_2 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M18 RDECO_2 RI_2 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M17 RDECO_1 RI_2 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M16 RDECO_0 RI_2 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M15 RDECO_7 RIB_1 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M14 RDECO_6 RIB_1 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M13 RDECO_3 RIB_1 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M12 RDECO_2 RIB_1 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M11 RDECO_5 RI_1 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M10 RDECO_4 RI_1 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M9 RDECO_1 RI_1 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M7 RDECO_7 RIB_0 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M6 RDECO_5 RIB_0 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M5 RDECO_3 RIB_0 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M4 RDECO_1 RIB_0 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M3 RDECO_6 RI_0 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M2 RDECO_4 RI_0 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1 RDECO_2 RI_0 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M0 RDECO_0 RI_0 0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS RDEC3TO8A_G4 
* FILE NAME: SRAM2_MUX_DEMUX_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: MUX_DEMUX.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:33 2007.
   
* TERMINAL MAPPING: BIT<0> = BIT_0
*                   BIT<1> = BIT_1
*                   BIT<2> = BIT_2
*                   BIT<3> = BIT_3
*                   BIT<4> = BIT_4
*                   BIT<5> = BIT_5
*                   BIT<6> = BIT_6
*                   BIT<7> = BIT_7
*                   BIT<8> = BIT_8
*                   BIT<9> = BIT_9
*                   BIT<10> = BIT_10
*                   BIT<11> = BIT_11
*                   BIT<12> = BIT_12
*                   BIT<13> = BIT_13
*                   BIT<14> = BIT_14
*                   BIT<15> = BIT_15
*                   BIT<16> = BIT_16
*                   BIT<17> = BIT_17
*                   BIT<18> = BIT_18
*                   BIT<19> = BIT_19
*                   BIT<20> = BIT_20
*                   BIT<21> = BIT_21
*                   BIT<22> = BIT_22
*                   BIT<23> = BIT_23
*                   BIT<24> = BIT_24
*                   BIT<25> = BIT_25
*                   BIT<26> = BIT_26
*                   BIT<27> = BIT_27
*                   BIT<28> = BIT_28
*                   BIT<29> = BIT_29
*                   BIT<30> = BIT_30
*                   BIT<31> = BIT_31
*                   BIT_B<0> = BIT_B_0
*                   BIT_B<1> = BIT_B_1
*                   BIT_B<2> = BIT_B_2
*                   BIT_B<3> = BIT_B_3
*                   BIT_B<4> = BIT_B_4
*                   BIT_B<5> = BIT_B_5
*                   BIT_B<6> = BIT_B_6
*                   BIT_B<7> = BIT_B_7
*                   BIT_B<8> = BIT_B_8
*                   BIT_B<9> = BIT_B_9
*                   BIT_B<10> = BIT_B_10
*                   BIT_B<11> = BIT_B_11
*                   BIT_B<12> = BIT_B_12
*                   BIT_B<13> = BIT_B_13
*                   BIT_B<14> = BIT_B_14
*                   BIT_B<15> = BIT_B_15
*                   BIT_B<16> = BIT_B_16
*                   BIT_B<17> = BIT_B_17
*                   BIT_B<18> = BIT_B_18
*                   BIT_B<19> = BIT_B_19
*                   BIT_B<20> = BIT_B_20
*                   BIT_B<21> = BIT_B_21
*                   BIT_B<22> = BIT_B_22
*                   BIT_B<23> = BIT_B_23
*                   BIT_B<24> = BIT_B_24
*                   BIT_B<25> = BIT_B_25
*                   BIT_B<26> = BIT_B_26
*                   BIT_B<27> = BIT_B_27
*                   BIT_B<28> = BIT_B_28
*                   BIT_B<29> = BIT_B_29
*                   BIT_B<30> = BIT_B_30
*                   BIT_B<31> = BIT_B_31
*                   BIT_B_LOWER<0> = BIT_B_LOWER_0
*                   BIT_B_LOWER<1> = BIT_B_LOWER_1
*                   BIT_B_LOWER<2> = BIT_B_LOWER_2
*                   BIT_B_LOWER<3> = BIT_B_LOWER_3
*                   BIT_B_LOWER<4> = BIT_B_LOWER_4
*                   BIT_B_LOWER<5> = BIT_B_LOWER_5
*                   BIT_B_LOWER<6> = BIT_B_LOWER_6
*                   BIT_B_LOWER<7> = BIT_B_LOWER_7
*                   BIT_B_LOWER<8> = BIT_B_LOWER_8
*                   BIT_B_LOWER<9> = BIT_B_LOWER_9
*                   BIT_B_LOWER<10> = BIT_B_LOWER_10
*                   BIT_B_LOWER<11> = BIT_B_LOWER_11
*                   BIT_B_LOWER<12> = BIT_B_LOWER_12
*                   BIT_B_LOWER<13> = BIT_B_LOWER_13
*                   BIT_B_LOWER<14> = BIT_B_LOWER_14
*                   BIT_B_LOWER<15> = BIT_B_LOWER_15
*                   BIT_B_LOWER<16> = BIT_B_LOWER_16
*                   BIT_B_LOWER<17> = BIT_B_LOWER_17
*                   BIT_B_LOWER<18> = BIT_B_LOWER_18
*                   BIT_B_LOWER<19> = BIT_B_LOWER_19
*                   BIT_B_LOWER<20> = BIT_B_LOWER_20
*                   BIT_B_LOWER<21> = BIT_B_LOWER_21
*                   BIT_B_LOWER<22> = BIT_B_LOWER_22
*                   BIT_B_LOWER<23> = BIT_B_LOWER_23
*                   BIT_B_LOWER<24> = BIT_B_LOWER_24
*                   BIT_B_LOWER<25> = BIT_B_LOWER_25
*                   BIT_B_LOWER<26> = BIT_B_LOWER_26
*                   BIT_B_LOWER<27> = BIT_B_LOWER_27
*                   BIT_B_LOWER<28> = BIT_B_LOWER_28
*                   BIT_B_LOWER<29> = BIT_B_LOWER_29
*                   BIT_B_LOWER<30> = BIT_B_LOWER_30
*                   BIT_B_LOWER<31> = BIT_B_LOWER_31
*                   BIT_LOWER<0> = BIT_LOWER_0
*                   BIT_LOWER<1> = BIT_LOWER_1
*                   BIT_LOWER<2> = BIT_LOWER_2
*                   BIT_LOWER<3> = BIT_LOWER_3
*                   BIT_LOWER<4> = BIT_LOWER_4
*                   BIT_LOWER<5> = BIT_LOWER_5
*                   BIT_LOWER<6> = BIT_LOWER_6
*                   BIT_LOWER<7> = BIT_LOWER_7
*                   BIT_LOWER<8> = BIT_LOWER_8
*                   BIT_LOWER<9> = BIT_LOWER_9
*                   BIT_LOWER<10> = BIT_LOWER_10
*                   BIT_LOWER<11> = BIT_LOWER_11
*                   BIT_LOWER<12> = BIT_LOWER_12
*                   BIT_LOWER<13> = BIT_LOWER_13
*                   BIT_LOWER<14> = BIT_LOWER_14
*                   BIT_LOWER<15> = BIT_LOWER_15
*                   BIT_LOWER<16> = BIT_LOWER_16
*                   BIT_LOWER<17> = BIT_LOWER_17
*                   BIT_LOWER<18> = BIT_LOWER_18
*                   BIT_LOWER<19> = BIT_LOWER_19
*                   BIT_LOWER<20> = BIT_LOWER_20
*                   BIT_LOWER<21> = BIT_LOWER_21
*                   BIT_LOWER<22> = BIT_LOWER_22
*                   BIT_LOWER<23> = BIT_LOWER_23
*                   BIT_LOWER<24> = BIT_LOWER_24
*                   BIT_LOWER<25> = BIT_LOWER_25
*                   BIT_LOWER<26> = BIT_LOWER_26
*                   BIT_LOWER<27> = BIT_LOWER_27
*                   BIT_LOWER<28> = BIT_LOWER_28
*                   BIT_LOWER<29> = BIT_LOWER_29
*                   BIT_LOWER<30> = BIT_LOWER_30
*                   BIT_LOWER<31> = BIT_LOWER_31
*                   COL = COL
.SUBCKT MUX_DEMUX_G17 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 BIT_8 
+BIT_9 BIT_10 BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 BIT_19 
+BIT_20 BIT_21 BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 BIT_30 
+BIT_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 
+BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 
+BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 
+BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 BIT_B_29 BIT_B_30 BIT_B_31 BIT_B_LOWER_0 
+BIT_B_LOWER_1 BIT_B_LOWER_2 BIT_B_LOWER_3 BIT_B_LOWER_4 BIT_B_LOWER_5 
+BIT_B_LOWER_6 BIT_B_LOWER_7 BIT_B_LOWER_8 BIT_B_LOWER_9 BIT_B_LOWER_10 
+BIT_B_LOWER_11 BIT_B_LOWER_12 BIT_B_LOWER_13 BIT_B_LOWER_14 BIT_B_LOWER_15 
+BIT_B_LOWER_16 BIT_B_LOWER_17 BIT_B_LOWER_18 BIT_B_LOWER_19 BIT_B_LOWER_20 
+BIT_B_LOWER_21 BIT_B_LOWER_22 BIT_B_LOWER_23 BIT_B_LOWER_24 BIT_B_LOWER_25 
+BIT_B_LOWER_26 BIT_B_LOWER_27 BIT_B_LOWER_28 BIT_B_LOWER_29 BIT_B_LOWER_30 
+BIT_B_LOWER_31 BIT_LOWER_0 BIT_LOWER_1 BIT_LOWER_2 BIT_LOWER_3 BIT_LOWER_4 
+BIT_LOWER_5 BIT_LOWER_6 BIT_LOWER_7 BIT_LOWER_8 BIT_LOWER_9 BIT_LOWER_10 
+BIT_LOWER_11 BIT_LOWER_12 BIT_LOWER_13 BIT_LOWER_14 BIT_LOWER_15 BIT_LOWER_16 
+BIT_LOWER_17 BIT_LOWER_18 BIT_LOWER_19 BIT_LOWER_20 BIT_LOWER_21 BIT_LOWER_22 
+BIT_LOWER_23 BIT_LOWER_24 BIT_LOWER_25 BIT_LOWER_26 BIT_LOWER_27 BIT_LOWER_28 
+BIT_LOWER_29 BIT_LOWER_30 BIT_LOWER_31 COL 
XI256 COL NET60 INV_1 
M1016 BIT_B_LOWER_27 NET60 BIT_B_27 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1017 BIT_B_LOWER_26 NET60 BIT_B_26 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1018 BIT_B_LOWER_25 NET60 BIT_B_25 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1019 BIT_B_LOWER_24 NET60 BIT_B_24 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1020 BIT_B_LOWER_23 NET60 BIT_B_23 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1021 BIT_B_LOWER_22 NET60 BIT_B_22 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1022 BIT_B_LOWER_21 NET60 BIT_B_21 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1023 BIT_B_LOWER_20 NET60 BIT_B_20 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1040 BIT_B_LOWER_3 NET60 BIT_B_3 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1041 BIT_B_LOWER_2 NET60 BIT_B_2 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1042 BIT_B_LOWER_1 NET60 BIT_B_1 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1043 BIT_B_LOWER_0 NET60 BIT_B_0 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1027 BIT_B_LOWER_16 NET60 BIT_B_16 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1026 BIT_B_LOWER_17 NET60 BIT_B_17 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1025 BIT_B_LOWER_18 NET60 BIT_B_18 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1024 BIT_B_LOWER_19 NET60 BIT_B_19 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1039 BIT_B_LOWER_4 NET60 BIT_B_4 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1031 BIT_B_LOWER_12 NET60 BIT_B_12 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1015 BIT_B_LOWER_28 NET60 BIT_B_28 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1014 BIT_B_LOWER_29 NET60 BIT_B_29 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1038 BIT_B_LOWER_5 NET60 BIT_B_5 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1013 BIT_B_LOWER_30 NET60 BIT_B_30 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1037 BIT_B_LOWER_6 NET60 BIT_B_6 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1030 BIT_B_LOWER_13 NET60 BIT_B_13 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1012 BIT_B_LOWER_31 NET60 BIT_B_31 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1036 BIT_B_LOWER_7 NET60 BIT_B_7 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1035 BIT_B_LOWER_8 NET60 BIT_B_8 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1029 BIT_B_LOWER_14 NET60 BIT_B_14 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1034 BIT_B_LOWER_9 NET60 BIT_B_9 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M534 BIT_LOWER_1 NET60 BIT_1 VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M535 BIT_LOWER_2 NET60 BIT_2 VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M536 BIT_LOWER_3 NET60 BIT_3 VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M537 BIT_LOWER_4 NET60 BIT_4 VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M538 BIT_LOWER_5 NET60 BIT_5 VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M539 BIT_LOWER_6 NET60 BIT_6 VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M540 BIT_LOWER_7 NET60 BIT_7 VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M541 BIT_LOWER_8 NET60 BIT_8 VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M542 BIT_LOWER_9 NET60 BIT_9 VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M543 BIT_LOWER_10 NET60 BIT_10 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M544 BIT_LOWER_11 NET60 BIT_11 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M545 BIT_LOWER_12 NET60 BIT_12 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M546 BIT_LOWER_13 NET60 BIT_13 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M547 BIT_LOWER_14 NET60 BIT_14 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M548 BIT_LOWER_15 NET60 BIT_15 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M549 BIT_LOWER_16 NET60 BIT_16 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M550 BIT_LOWER_17 NET60 BIT_17 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M551 BIT_LOWER_18 NET60 BIT_18 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M552 BIT_LOWER_19 NET60 BIT_19 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M553 BIT_LOWER_20 NET60 BIT_20 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M554 BIT_LOWER_21 NET60 BIT_21 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M555 BIT_LOWER_22 NET60 BIT_22 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M556 BIT_LOWER_23 NET60 BIT_23 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M557 BIT_LOWER_24 NET60 BIT_24 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M558 BIT_LOWER_25 NET60 BIT_25 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M559 BIT_LOWER_26 NET60 BIT_26 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M560 BIT_LOWER_27 NET60 BIT_27 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M561 BIT_LOWER_28 NET60 BIT_28 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M562 BIT_LOWER_29 NET60 BIT_29 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M563 BIT_LOWER_30 NET60 BIT_30 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M564 BIT_LOWER_31 NET60 BIT_31 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1032 BIT_B_LOWER_11 NET60 BIT_B_11 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1028 BIT_B_LOWER_15 NET60 BIT_B_15 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1033 BIT_B_LOWER_10 NET60 BIT_B_10 VDD!  PFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1 BIT_LOWER_0 NET60 BIT_0 VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1291 BIT_B_8 COL BIT_B_LOWER_8 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1292 BIT_B_7 COL BIT_B_LOWER_7 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1293 BIT_B_6 COL BIT_B_LOWER_6 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1294 BIT_B_5 COL BIT_B_LOWER_5 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1295 BIT_B_4 COL BIT_B_LOWER_4 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1296 BIT_B_3 COL BIT_B_LOWER_3 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1297 BIT_B_2 COL BIT_B_LOWER_2 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1298 BIT_B_1 COL BIT_B_LOWER_1 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1299 BIT_B_0 COL BIT_B_LOWER_0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1290 BIT_B_9 COL BIT_B_LOWER_9 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1289 BIT_B_10 COL BIT_B_LOWER_10 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1274 BIT_B_25 COL BIT_B_LOWER_25 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1288 BIT_B_11 COL BIT_B_LOWER_11 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1287 BIT_B_12 COL BIT_B_LOWER_12 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1273 BIT_B_26 COL BIT_B_LOWER_26 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1286 BIT_B_13 COL BIT_B_LOWER_13 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1285 BIT_B_14 COL BIT_B_LOWER_14 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1272 BIT_B_27 COL BIT_B_LOWER_27 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1284 BIT_B_15 COL BIT_B_LOWER_15 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1283 BIT_B_16 COL BIT_B_LOWER_16 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1271 BIT_B_28 COL BIT_B_LOWER_28 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1282 BIT_B_17 COL BIT_B_LOWER_17 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1281 BIT_B_18 COL BIT_B_LOWER_18 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1270 BIT_B_29 COL BIT_B_LOWER_29 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1280 BIT_B_19 COL BIT_B_LOWER_19 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1279 BIT_B_20 COL BIT_B_LOWER_20 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1269 BIT_B_30 COL BIT_B_LOWER_30 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M502 BIT_1 COL BIT_LOWER_1 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M503 BIT_2 COL BIT_LOWER_2 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M504 BIT_3 COL BIT_LOWER_3 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M505 BIT_4 COL BIT_LOWER_4 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M506 BIT_5 COL BIT_LOWER_5 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M507 BIT_6 COL BIT_LOWER_6 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M508 BIT_7 COL BIT_LOWER_7 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M509 BIT_8 COL BIT_LOWER_8 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M510 BIT_9 COL BIT_LOWER_9 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M511 BIT_10 COL BIT_LOWER_10 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M512 BIT_11 COL BIT_LOWER_11 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M513 BIT_12 COL BIT_LOWER_12 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M514 BIT_13 COL BIT_LOWER_13 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M515 BIT_14 COL BIT_LOWER_14 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M516 BIT_15 COL BIT_LOWER_15 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M517 BIT_16 COL BIT_LOWER_16 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M518 BIT_17 COL BIT_LOWER_17 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M519 BIT_18 COL BIT_LOWER_18 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M520 BIT_19 COL BIT_LOWER_19 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M521 BIT_20 COL BIT_LOWER_20 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M522 BIT_21 COL BIT_LOWER_21 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M523 BIT_22 COL BIT_LOWER_22 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M524 BIT_23 COL BIT_LOWER_23 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M525 BIT_24 COL BIT_LOWER_24 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M526 BIT_25 COL BIT_LOWER_25 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M527 BIT_26 COL BIT_LOWER_26 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M528 BIT_27 COL BIT_LOWER_27 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M529 BIT_28 COL BIT_LOWER_28 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M530 BIT_29 COL BIT_LOWER_29 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M531 BIT_30 COL BIT_LOWER_30 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M532 BIT_31 COL BIT_LOWER_31 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M1275 BIT_B_24 COL BIT_B_LOWER_24 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1276 BIT_B_23 COL BIT_B_LOWER_23 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1268 BIT_B_31 COL BIT_B_LOWER_31 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1277 BIT_B_22 COL BIT_B_LOWER_22 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M1278 BIT_B_21 COL BIT_B_LOWER_21 0  NFET  L=200E-9 W=400E-9 
+AD=+2.00000000E-13 AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 
+NRD=+1.25000000E+00 NRS=+1.25000000E+00 M=1.0 
M0 BIT_0 COL BIT_LOWER_0 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
   
   
* FILE NAME: SRAM2_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_1 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(4E-6) AD=+2.00000000E-12 
+AS=+2.00000000E-12 PD=+9.00000000E-06 PS=+9.00000000E-06 NRD=+1.25000000E-01 
+NRS=+1.25000000E-01 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(2E-6) AD=+1.00000000E-12 AS=+1.00000000E-12 
+PD=+5.00000000E-06 PS=+5.00000000E-06 NRD=+2.50000000E-01 NRS=+2.50000000E-01 
+M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS MUX_DEMUX_G17 
* FILE NAME: SRAM_RDEC6TO64_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: RDEC6TO64.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:39 2007.
   
* TERMINAL MAPPING: RDECO<0> = RDECO_0
*                   RDECO<1> = RDECO_1
*                   RDECO<2> = RDECO_2
*                   RDECO<3> = RDECO_3
*                   RDECO<4> = RDECO_4
*                   RDECO<5> = RDECO_5
*                   RDECO<6> = RDECO_6
*                   RDECO<7> = RDECO_7
*                   RDECO<8> = RDECO_8
*                   RDECO<9> = RDECO_9
*                   RDECO<10> = RDECO_10
*                   RDECO<11> = RDECO_11
*                   RDECO<12> = RDECO_12
*                   RDECO<13> = RDECO_13
*                   RDECO<14> = RDECO_14
*                   RDECO<15> = RDECO_15
*                   RDECO<16> = RDECO_16
*                   RDECO<17> = RDECO_17
*                   RDECO<18> = RDECO_18
*                   RDECO<19> = RDECO_19
*                   RDECO<20> = RDECO_20
*                   RDECO<21> = RDECO_21
*                   RDECO<22> = RDECO_22
*                   RDECO<23> = RDECO_23
*                   RDECO<24> = RDECO_24
*                   RDECO<25> = RDECO_25
*                   RDECO<26> = RDECO_26
*                   RDECO<27> = RDECO_27
*                   RDECO<28> = RDECO_28
*                   RDECO<29> = RDECO_29
*                   RDECO<30> = RDECO_30
*                   RDECO<31> = RDECO_31
*                   RDECO<32> = RDECO_32
*                   RDECO<33> = RDECO_33
*                   RDECO<34> = RDECO_34
*                   RDECO<35> = RDECO_35
*                   RDECO<36> = RDECO_36
*                   RDECO<37> = RDECO_37
*                   RDECO<38> = RDECO_38
*                   RDECO<39> = RDECO_39
*                   RDECO<40> = RDECO_40
*                   RDECO<41> = RDECO_41
*                   RDECO<42> = RDECO_42
*                   RDECO<43> = RDECO_43
*                   RDECO<44> = RDECO_44
*                   RDECO<45> = RDECO_45
*                   RDECO<46> = RDECO_46
*                   RDECO<47> = RDECO_47
*                   RDECO<48> = RDECO_48
*                   RDECO<49> = RDECO_49
*                   RDECO<50> = RDECO_50
*                   RDECO<51> = RDECO_51
*                   RDECO<52> = RDECO_52
*                   RDECO<53> = RDECO_53
*                   RDECO<54> = RDECO_54
*                   RDECO<55> = RDECO_55
*                   RDECO<56> = RDECO_56
*                   RDECO<57> = RDECO_57
*                   RDECO<58> = RDECO_58
*                   RDECO<59> = RDECO_59
*                   RDECO<60> = RDECO_60
*                   RDECO<61> = RDECO_61
*                   RDECO<62> = RDECO_62
*                   RDECO<63> = RDECO_63
*                   RI<0> = RI_0
*                   RI<1> = RI_1
*                   RI<2> = RI_2
*                   RI<3> = RI_3
*                   RI<4> = RI_4
*                   RI<5> = RI_5
*                   RIB<0> = RIB_0
*                   RIB<1> = RIB_1
*                   RIB<2> = RIB_2
*                   RIB<3> = RIB_3
*                   RIB<4> = RIB_4
*                   RIB<5> = RIB_5
*                   TOP = TOP
.SUBCKT RDEC6TO64_G10 RDECO_0 RDECO_1 RDECO_2 RDECO_3 RDECO_4 RDECO_5 RDECO_6 
+RDECO_7 RDECO_8 RDECO_9 RDECO_10 RDECO_11 RDECO_12 RDECO_13 RDECO_14 RDECO_15 
+RDECO_16 RDECO_17 RDECO_18 RDECO_19 RDECO_20 RDECO_21 RDECO_22 RDECO_23 
+RDECO_24 RDECO_25 RDECO_26 RDECO_27 RDECO_28 RDECO_29 RDECO_30 RDECO_31 
+RDECO_32 RDECO_33 RDECO_34 RDECO_35 RDECO_36 RDECO_37 RDECO_38 RDECO_39 
+RDECO_40 RDECO_41 RDECO_42 RDECO_43 RDECO_44 RDECO_45 RDECO_46 RDECO_47 
+RDECO_48 RDECO_49 RDECO_50 RDECO_51 RDECO_52 RDECO_53 RDECO_54 RDECO_55 
+RDECO_56 RDECO_57 RDECO_58 RDECO_59 RDECO_60 RDECO_61 RDECO_62 RDECO_63 RI_0 
+RI_1 RI_2 RI_3 RI_4 RI_5 RIB_0 RIB_1 RIB_2 RIB_3 RIB_4 RIB_5 TOP 
M66 RDECO_63 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M67 RDECO_62 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M68 RDECO_61 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M69 RDECO_60 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M70 RDECO_59 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M71 RDECO_58 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M72 RDECO_57 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M73 RDECO_56 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M74 RDECO_55 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M75 RDECO_54 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M76 RDECO_53 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M77 RDECO_52 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M78 RDECO_51 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M79 RDECO_50 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M80 RDECO_49 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M81 RDECO_48 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M82 RDECO_47 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M83 RDECO_46 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M84 RDECO_45 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M85 RDECO_44 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M86 RDECO_43 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M87 RDECO_42 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M88 RDECO_41 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M89 RDECO_40 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M90 RDECO_39 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M91 RDECO_38 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M92 RDECO_37 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M93 RDECO_36 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M94 RDECO_35 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M95 RDECO_34 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M96 RDECO_32 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M97 RDECO_33 RIB_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M33 RDECO_31 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M32 RDECO_30 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M31 RDECO_29 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M30 RDECO_28 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M29 RDECO_27 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M28 RDECO_26 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M27 RDECO_25 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M26 RDECO_24 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M25 RDECO_23 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M24 RDECO_22 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M23 RDECO_21 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M22 RDECO_20 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M21 RDECO_19 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M20 RDECO_18 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M19 RDECO_17 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M18 RDECO_16 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M17 RDECO_15 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M16 RDECO_14 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M15 RDECO_13 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M14 RDECO_12 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M7 RDECO_5 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M6 RDECO_4 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M5 RDECO_3 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M4 RDECO_2 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M3 RDECO_1 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M2 RDECO_0 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M8 RDECO_6 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M10 RDECO_8 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M9 RDECO_7 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M12 RDECO_10 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M11 RDECO_9 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M13 RDECO_11 RI_5 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
XI12 RDECO_32 RDECO_33 RDECO_34 RDECO_35 RDECO_36 RDECO_37 RDECO_38 RDECO_39 
+RDECO_40 RDECO_41 RDECO_42 RDECO_43 RDECO_44 RDECO_45 RDECO_46 RDECO_47 
+RDECO_48 RDECO_49 RDECO_50 RDECO_51 RDECO_52 RDECO_53 RDECO_54 RDECO_55 
+RDECO_56 RDECO_57 RDECO_58 RDECO_59 RDECO_60 RDECO_61 RDECO_62 RDECO_63 RI_0 
+RI_1 RI_2 RI_3 RI_4 RIB_0 RIB_1 RIB_2 RIB_3 RIB_4 NET76 RDEC5TO32_G9 
XI11 RDECO_0 RDECO_1 RDECO_2 RDECO_3 RDECO_4 RDECO_5 RDECO_6 RDECO_7 RDECO_8 
+RDECO_9 RDECO_10 RDECO_11 RDECO_12 RDECO_13 RDECO_14 RDECO_15 RDECO_16 
+RDECO_17 RDECO_18 RDECO_19 RDECO_20 RDECO_21 RDECO_22 RDECO_23 RDECO_24 
+RDECO_25 RDECO_26 RDECO_27 RDECO_28 RDECO_29 RDECO_30 RDECO_31 RI_0 RI_1 RI_2 
+RI_3 RI_4 RIB_0 RIB_1 RIB_2 RIB_3 RIB_4 NET33 RDEC5TO32_G9 
M1 NET76 RIB_5 TOP VDD!  PFET  L=200E-9 W=147.2E-6 AD=+7.36000000E-11 
+AS=+7.36000000E-11 PD=+2.95400000E-04 PS=+2.95400000E-04 NRD=+3.39673913E-03 
+NRS=+3.39673913E-03 M=1.0 
M0 NET33 RI_5 TOP VDD!  PFET  L=200E-9 W=147.2E-6 AD=+7.36000000E-11 
+AS=+7.36000000E-11 PD=+2.95400000E-04 PS=+2.95400000E-04 NRD=+3.39673913E-03 
+NRS=+3.39673913E-03 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS RDEC6TO64_G10 
* FILE NAME: SRAM2_T1_PI_MODEL64_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: T1_PI_MODEL64.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:36 2007.
   
* TERMINAL MAPPING: IN<0> = IN_0
*                   IN<1> = IN_1
*                   IN<2> = IN_2
*                   IN<3> = IN_3
*                   IN<4> = IN_4
*                   IN<5> = IN_5
*                   IN<6> = IN_6
*                   IN<7> = IN_7
*                   IN<8> = IN_8
*                   IN<9> = IN_9
*                   IN<10> = IN_10
*                   IN<11> = IN_11
*                   IN<12> = IN_12
*                   IN<13> = IN_13
*                   IN<14> = IN_14
*                   IN<15> = IN_15
*                   IN<16> = IN_16
*                   IN<17> = IN_17
*                   IN<18> = IN_18
*                   IN<19> = IN_19
*                   IN<20> = IN_20
*                   IN<21> = IN_21
*                   IN<22> = IN_22
*                   IN<23> = IN_23
*                   IN<24> = IN_24
*                   IN<25> = IN_25
*                   IN<26> = IN_26
*                   IN<27> = IN_27
*                   IN<28> = IN_28
*                   IN<29> = IN_29
*                   IN<30> = IN_30
*                   IN<31> = IN_31
*                   IN<32> = IN_32
*                   IN<33> = IN_33
*                   IN<34> = IN_34
*                   IN<35> = IN_35
*                   IN<36> = IN_36
*                   IN<37> = IN_37
*                   IN<38> = IN_38
*                   IN<39> = IN_39
*                   IN<40> = IN_40
*                   IN<41> = IN_41
*                   IN<42> = IN_42
*                   IN<43> = IN_43
*                   IN<44> = IN_44
*                   IN<45> = IN_45
*                   IN<46> = IN_46
*                   IN<47> = IN_47
*                   IN<48> = IN_48
*                   IN<49> = IN_49
*                   IN<50> = IN_50
*                   IN<51> = IN_51
*                   IN<52> = IN_52
*                   IN<53> = IN_53
*                   IN<54> = IN_54
*                   IN<55> = IN_55
*                   IN<56> = IN_56
*                   IN<57> = IN_57
*                   IN<58> = IN_58
*                   IN<59> = IN_59
*                   IN<60> = IN_60
*                   IN<61> = IN_61
*                   IN<62> = IN_62
*                   IN<63> = IN_63
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
*                   OUT<3> = OUT_3
*                   OUT<4> = OUT_4
*                   OUT<5> = OUT_5
*                   OUT<6> = OUT_6
*                   OUT<7> = OUT_7
*                   OUT<8> = OUT_8
*                   OUT<9> = OUT_9
*                   OUT<10> = OUT_10
*                   OUT<11> = OUT_11
*                   OUT<12> = OUT_12
*                   OUT<13> = OUT_13
*                   OUT<14> = OUT_14
*                   OUT<15> = OUT_15
*                   OUT<16> = OUT_16
*                   OUT<17> = OUT_17
*                   OUT<18> = OUT_18
*                   OUT<19> = OUT_19
*                   OUT<20> = OUT_20
*                   OUT<21> = OUT_21
*                   OUT<22> = OUT_22
*                   OUT<23> = OUT_23
*                   OUT<24> = OUT_24
*                   OUT<25> = OUT_25
*                   OUT<26> = OUT_26
*                   OUT<27> = OUT_27
*                   OUT<28> = OUT_28
*                   OUT<29> = OUT_29
*                   OUT<30> = OUT_30
*                   OUT<31> = OUT_31
*                   OUT<32> = OUT_32
*                   OUT<33> = OUT_33
*                   OUT<34> = OUT_34
*                   OUT<35> = OUT_35
*                   OUT<36> = OUT_36
*                   OUT<37> = OUT_37
*                   OUT<38> = OUT_38
*                   OUT<39> = OUT_39
*                   OUT<40> = OUT_40
*                   OUT<41> = OUT_41
*                   OUT<42> = OUT_42
*                   OUT<43> = OUT_43
*                   OUT<44> = OUT_44
*                   OUT<45> = OUT_45
*                   OUT<46> = OUT_46
*                   OUT<47> = OUT_47
*                   OUT<48> = OUT_48
*                   OUT<49> = OUT_49
*                   OUT<50> = OUT_50
*                   OUT<51> = OUT_51
*                   OUT<52> = OUT_52
*                   OUT<53> = OUT_53
*                   OUT<54> = OUT_54
*                   OUT<55> = OUT_55
*                   OUT<56> = OUT_56
*                   OUT<57> = OUT_57
*                   OUT<58> = OUT_58
*                   OUT<59> = OUT_59
*                   OUT<60> = OUT_60
*                   OUT<61> = OUT_61
*                   OUT<62> = OUT_62
*                   OUT<63> = OUT_63
.SUBCKT SUB1 IN_0 IN_1 IN_2 IN_3 IN_4 IN_5 IN_6 IN_7 IN_8 IN_9 IN_10 IN_11 
+IN_12 IN_13 IN_14 IN_15 IN_16 IN_17 IN_18 IN_19 IN_20 IN_21 IN_22 IN_23 IN_24 
+IN_25 IN_26 IN_27 IN_28 IN_29 IN_30 IN_31 IN_32 IN_33 IN_34 IN_35 IN_36 IN_37 
+IN_38 IN_39 IN_40 IN_41 IN_42 IN_43 IN_44 IN_45 IN_46 IN_47 IN_48 IN_49 IN_50 
+IN_51 IN_52 IN_53 IN_54 IN_55 IN_56 IN_57 IN_58 IN_59 IN_60 IN_61 IN_62 IN_63 
+OUT_0 OUT_1 OUT_2 OUT_3 OUT_4 OUT_5 OUT_6 OUT_7 OUT_8 OUT_9 OUT_10 OUT_11 
+OUT_12 OUT_13 OUT_14 OUT_15 OUT_16 OUT_17 OUT_18 OUT_19 OUT_20 OUT_21 OUT_22 
+OUT_23 OUT_24 OUT_25 OUT_26 OUT_27 OUT_28 OUT_29 OUT_30 OUT_31 OUT_32 OUT_33 
+OUT_34 OUT_35 OUT_36 OUT_37 OUT_38 OUT_39 OUT_40 OUT_41 OUT_42 OUT_43 OUT_44 
+OUT_45 OUT_46 OUT_47 OUT_48 OUT_49 OUT_50 OUT_51 OUT_52 OUT_53 OUT_54 OUT_55 
+OUT_56 OUT_57 OUT_58 OUT_59 OUT_60 OUT_61 OUT_62 OUT_63 
XI32 IN_32 OUT_32 TL_PI_MODEL_1 
XI33 IN_33 OUT_33 TL_PI_MODEL_1 
XI34 IN_34 OUT_34 TL_PI_MODEL_1 
XI35 IN_35 OUT_35 TL_PI_MODEL_1 
XI36 IN_36 OUT_36 TL_PI_MODEL_1 
XI37 IN_37 OUT_37 TL_PI_MODEL_1 
XI38 IN_38 OUT_38 TL_PI_MODEL_1 
XI39 IN_39 OUT_39 TL_PI_MODEL_1 
XI40 IN_40 OUT_40 TL_PI_MODEL_1 
XI41 IN_41 OUT_41 TL_PI_MODEL_1 
XI42 IN_42 OUT_42 TL_PI_MODEL_1 
XI43 IN_43 OUT_43 TL_PI_MODEL_1 
XI44 IN_44 OUT_44 TL_PI_MODEL_1 
XI45 IN_45 OUT_45 TL_PI_MODEL_1 
XI46 IN_46 OUT_46 TL_PI_MODEL_1 
XI47 IN_47 OUT_47 TL_PI_MODEL_1 
XI48 IN_48 OUT_48 TL_PI_MODEL_1 
XI49 IN_49 OUT_49 TL_PI_MODEL_1 
XI50 IN_50 OUT_50 TL_PI_MODEL_1 
XI51 IN_51 OUT_51 TL_PI_MODEL_1 
XI52 IN_52 OUT_52 TL_PI_MODEL_1 
XI53 IN_53 OUT_53 TL_PI_MODEL_1 
XI54 IN_54 OUT_54 TL_PI_MODEL_1 
XI55 IN_55 OUT_55 TL_PI_MODEL_1 
XI56 IN_56 OUT_56 TL_PI_MODEL_1 
XI57 IN_57 OUT_57 TL_PI_MODEL_1 
XI58 IN_58 OUT_58 TL_PI_MODEL_1 
XI59 IN_59 OUT_59 TL_PI_MODEL_1 
XI60 IN_60 OUT_60 TL_PI_MODEL_1 
XI61 IN_61 OUT_61 TL_PI_MODEL_1 
XI62 IN_62 OUT_62 TL_PI_MODEL_1 
XI63 IN_63 OUT_63 TL_PI_MODEL_1 
XI31 IN_31 OUT_31 TL_PI_MODEL_1 
XI30 IN_30 OUT_30 TL_PI_MODEL_1 
XI29 IN_29 OUT_29 TL_PI_MODEL_1 
XI28 IN_28 OUT_28 TL_PI_MODEL_1 
XI27 IN_27 OUT_27 TL_PI_MODEL_1 
XI26 IN_26 OUT_26 TL_PI_MODEL_1 
XI25 IN_25 OUT_25 TL_PI_MODEL_1 
XI24 IN_24 OUT_24 TL_PI_MODEL_1 
XI23 IN_23 OUT_23 TL_PI_MODEL_1 
XI22 IN_22 OUT_22 TL_PI_MODEL_1 
XI21 IN_21 OUT_21 TL_PI_MODEL_1 
XI20 IN_20 OUT_20 TL_PI_MODEL_1 
XI19 IN_19 OUT_19 TL_PI_MODEL_1 
XI18 IN_18 OUT_18 TL_PI_MODEL_1 
XI17 IN_17 OUT_17 TL_PI_MODEL_1 
XI16 IN_16 OUT_16 TL_PI_MODEL_1 
XI15 IN_15 OUT_15 TL_PI_MODEL_1 
XI14 IN_14 OUT_14 TL_PI_MODEL_1 
XI13 IN_13 OUT_13 TL_PI_MODEL_1 
XI12 IN_12 OUT_12 TL_PI_MODEL_1 
XI11 IN_11 OUT_11 TL_PI_MODEL_1 
XI10 IN_10 OUT_10 TL_PI_MODEL_1 
XI9 IN_9 OUT_9 TL_PI_MODEL_1 
XI8 IN_8 OUT_8 TL_PI_MODEL_1 
XI7 IN_7 OUT_7 TL_PI_MODEL_1 
XI6 IN_6 OUT_6 TL_PI_MODEL_1 
XI5 IN_5 OUT_5 TL_PI_MODEL_1 
XI4 IN_4 OUT_4 TL_PI_MODEL_1 
XI3 IN_3 OUT_3 TL_PI_MODEL_1 
XI2 IN_2 OUT_2 TL_PI_MODEL_1 
XI1 IN_1 OUT_1 TL_PI_MODEL_1 
XI0 IN_0 OUT_0 TL_PI_MODEL_1 
   
   
* FILE NAME: SRAM2_TL_PI_MODEL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:31 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT TL_PI_MODEL_1 IN OUT 
C0 IN 0  (291E-15) M=1.0 
C1 OUT 0  (291E-15) M=1.0 
R0 IN OUT  (204.8) M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SUB1 
* FILE NAME: SRAM2_CONTROL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: CONTROL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:35 2007.
   
* TERMINAL MAPPING: IN<0> = IN_0
*                   IN<1> = IN_1
*                   IN<2> = IN_2
*                   IN<3> = IN_3
*                   IN<4> = IN_4
*                   IN<5> = IN_5
*                   IN<6> = IN_6
*                   IN<7> = IN_7
*                   IN<8> = IN_8
*                   IN<9> = IN_9
*                   IN<10> = IN_10
*                   IN<11> = IN_11
*                   IN<12> = IN_12
*                   IN<13> = IN_13
*                   IN<14> = IN_14
*                   IN<15> = IN_15
*                   IN<16> = IN_16
*                   IN<17> = IN_17
*                   IN<18> = IN_18
*                   IN<19> = IN_19
*                   IN<20> = IN_20
*                   IN<21> = IN_21
*                   IN<22> = IN_22
*                   IN<23> = IN_23
*                   IN<24> = IN_24
*                   IN<25> = IN_25
*                   IN<26> = IN_26
*                   IN<27> = IN_27
*                   IN<28> = IN_28
*                   IN<29> = IN_29
*                   IN<30> = IN_30
*                   IN<31> = IN_31
*                   IN<32> = IN_32
*                   IN<33> = IN_33
*                   IN<34> = IN_34
*                   IN<35> = IN_35
*                   IN<36> = IN_36
*                   IN<37> = IN_37
*                   IN<38> = IN_38
*                   IN<39> = IN_39
*                   IN<40> = IN_40
*                   IN<41> = IN_41
*                   IN<42> = IN_42
*                   IN<43> = IN_43
*                   IN<44> = IN_44
*                   IN<45> = IN_45
*                   IN<46> = IN_46
*                   IN<47> = IN_47
*                   IN<48> = IN_48
*                   IN<49> = IN_49
*                   IN<50> = IN_50
*                   IN<51> = IN_51
*                   IN<52> = IN_52
*                   IN<53> = IN_53
*                   IN<54> = IN_54
*                   IN<55> = IN_55
*                   IN<56> = IN_56
*                   IN<57> = IN_57
*                   IN<58> = IN_58
*                   IN<59> = IN_59
*                   IN<60> = IN_60
*                   IN<61> = IN_61
*                   IN<62> = IN_62
*                   IN<63> = IN_63
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
*                   OUT<3> = OUT_3
*                   OUT<4> = OUT_4
*                   OUT<5> = OUT_5
*                   OUT<6> = OUT_6
*                   OUT<7> = OUT_7
*                   OUT<8> = OUT_8
*                   OUT<9> = OUT_9
*                   OUT<10> = OUT_10
*                   OUT<11> = OUT_11
*                   OUT<12> = OUT_12
*                   OUT<13> = OUT_13
*                   OUT<14> = OUT_14
*                   OUT<15> = OUT_15
*                   OUT<16> = OUT_16
*                   OUT<17> = OUT_17
*                   OUT<18> = OUT_18
*                   OUT<19> = OUT_19
*                   OUT<20> = OUT_20
*                   OUT<21> = OUT_21
*                   OUT<22> = OUT_22
*                   OUT<23> = OUT_23
*                   OUT<24> = OUT_24
*                   OUT<25> = OUT_25
*                   OUT<26> = OUT_26
*                   OUT<27> = OUT_27
*                   OUT<28> = OUT_28
*                   OUT<29> = OUT_29
*                   OUT<30> = OUT_30
*                   OUT<31> = OUT_31
*                   OUT<32> = OUT_32
*                   OUT<33> = OUT_33
*                   OUT<34> = OUT_34
*                   OUT<35> = OUT_35
*                   OUT<36> = OUT_36
*                   OUT<37> = OUT_37
*                   OUT<38> = OUT_38
*                   OUT<39> = OUT_39
*                   OUT<40> = OUT_40
*                   OUT<41> = OUT_41
*                   OUT<42> = OUT_42
*                   OUT<43> = OUT_43
*                   OUT<44> = OUT_44
*                   OUT<45> = OUT_45
*                   OUT<46> = OUT_46
*                   OUT<47> = OUT_47
*                   OUT<48> = OUT_48
*                   OUT<49> = OUT_49
*                   OUT<50> = OUT_50
*                   OUT<51> = OUT_51
*                   OUT<52> = OUT_52
*                   OUT<53> = OUT_53
*                   OUT<54> = OUT_54
*                   OUT<55> = OUT_55
*                   OUT<56> = OUT_56
*                   OUT<57> = OUT_57
*                   OUT<58> = OUT_58
*                   OUT<59> = OUT_59
*                   OUT<60> = OUT_60
*                   OUT<61> = OUT_61
*                   OUT<62> = OUT_62
*                   OUT<63> = OUT_63
*                   WORD_EN = WORD_EN
.SUBCKT CONTROL_G19 IN_0 IN_1 IN_2 IN_3 IN_4 IN_5 IN_6 IN_7 IN_8 IN_9 IN_10 
+IN_11 IN_12 IN_13 IN_14 IN_15 IN_16 IN_17 IN_18 IN_19 IN_20 IN_21 IN_22 IN_23 
+IN_24 IN_25 IN_26 IN_27 IN_28 IN_29 IN_30 IN_31 IN_32 IN_33 IN_34 IN_35 IN_36 
+IN_37 IN_38 IN_39 IN_40 IN_41 IN_42 IN_43 IN_44 IN_45 IN_46 IN_47 IN_48 IN_49 
+IN_50 IN_51 IN_52 IN_53 IN_54 IN_55 IN_56 IN_57 IN_58 IN_59 IN_60 IN_61 IN_62 
+IN_63 OUT_0 OUT_1 OUT_2 OUT_3 OUT_4 OUT_5 OUT_6 OUT_7 OUT_8 OUT_9 OUT_10 
+OUT_11 OUT_12 OUT_13 OUT_14 OUT_15 OUT_16 OUT_17 OUT_18 OUT_19 OUT_20 OUT_21 
+OUT_22 OUT_23 OUT_24 OUT_25 OUT_26 OUT_27 OUT_28 OUT_29 OUT_30 OUT_31 OUT_32 
+OUT_33 OUT_34 OUT_35 OUT_36 OUT_37 OUT_38 OUT_39 OUT_40 OUT_41 OUT_42 OUT_43 
+OUT_44 OUT_45 OUT_46 OUT_47 OUT_48 OUT_49 OUT_50 OUT_51 OUT_52 OUT_53 OUT_54 
+OUT_55 OUT_56 OUT_57 OUT_58 OUT_59 OUT_60 OUT_61 OUT_62 OUT_63 WORD_EN 
XI449 NET0363 OUT_49 INV_1 
XI453 NET0357 OUT_50 INV_1 
XI457 NET0697 OUT_51 INV_1 
XI461 NET0345 OUT_52 INV_1 
XI465 NET0691 OUT_53 INV_1 
XI469 NET0333 OUT_54 INV_1 
XI473 NET0685 OUT_55 INV_1 
XI477 NET0682 OUT_56 INV_1 
XI481 NET0679 OUT_57 INV_1 
XI485 NET0676 OUT_58 INV_1 
XI489 NET0303 OUT_59 INV_1 
XI493 NET0297 OUT_60 INV_1 
XI497 NET0291 OUT_61 INV_1 
XI501 NET0285 OUT_62 INV_1 
XI505 NET0279 OUT_63 INV_1 
XI257 NET0847 OUT_1 INV_1 
XI261 NET0645 OUT_2 INV_1 
XI289 NET0603 OUT_9 INV_1 
XI441 NET0709 OUT_47 INV_1 
XI437 NET0712 OUT_46 INV_1 
XI269 NET0633 OUT_4 INV_1 
XI301 NET0585 OUT_12 INV_1 
XI365 NET0766 OUT_28 INV_1 
XI445 NET0369 OUT_48 INV_1 
XI277 NET0621 OUT_6 INV_1 
XI273 NET0627 OUT_5 INV_1 
XI281 NET0829 OUT_7 INV_1 
XI285 NET0826 OUT_8 INV_1 
XI309 NET0573 OUT_14 INV_1 
XI313 NET0805 OUT_15 INV_1 
XI265 NET0841 OUT_3 INV_1 
XI293 NET0597 OUT_10 INV_1 
XI305 NET0579 OUT_13 INV_1 
XI433 NET0715 OUT_45 INV_1 
XI373 NET0760 OUT_30 INV_1 
XI317 NET0561 OUT_16 INV_1 
XI377 NET0757 OUT_31 INV_1 
XI321 NET0555 OUT_17 INV_1 
XI381 NET0754 OUT_32 INV_1 
XI325 NET0549 OUT_18 INV_1 
XI385 NET0459 OUT_33 INV_1 
XI329 NET0543 OUT_19 INV_1 
XI389 NET0453 OUT_34 INV_1 
XI333 NET0537 OUT_20 INV_1 
XI393 NET0745 OUT_35 INV_1 
XI337 NET0531 OUT_21 INV_1 
XI397 NET0742 OUT_36 INV_1 
XI341 NET0525 OUT_22 INV_1 
XI401 NET0435 OUT_37 INV_1 
XI345 NET0519 OUT_23 INV_1 
XI405 NET0429 OUT_38 INV_1 
XI349 NET0778 OUT_24 INV_1 
XI409 NET0733 OUT_39 INV_1 
XI353 NET0775 OUT_25 INV_1 
XI413 NET0417 OUT_40 INV_1 
XI357 NET0501 OUT_26 INV_1 
XI417 NET0727 OUT_41 INV_1 
XI361 NET0495 OUT_27 INV_1 
XI297 NET0817 OUT_11 INV_1 
XI421 NET0405 OUT_42 INV_1 
XI425 NET0399 OUT_43 INV_1 
XI369 NET0763 OUT_29 INV_1 
XI429 NET0718 OUT_44 INV_1 
XI1 NET50 OUT_0 INV_1 
XI448 WORD_EN IN_49 NET0363 NAND2_2 
XI452 WORD_EN IN_50 NET0357 NAND2_2 
XI456 WORD_EN IN_51 NET0697 NAND2_2 
XI460 WORD_EN IN_52 NET0345 NAND2_2 
XI464 WORD_EN IN_53 NET0691 NAND2_2 
XI468 WORD_EN IN_54 NET0333 NAND2_2 
XI472 WORD_EN IN_55 NET0685 NAND2_2 
XI476 WORD_EN IN_56 NET0682 NAND2_2 
XI480 WORD_EN IN_57 NET0679 NAND2_2 
XI484 WORD_EN IN_58 NET0676 NAND2_2 
XI488 WORD_EN IN_59 NET0303 NAND2_2 
XI492 WORD_EN IN_60 NET0297 NAND2_2 
XI496 WORD_EN IN_61 NET0291 NAND2_2 
XI500 WORD_EN IN_62 NET0285 NAND2_2 
XI504 WORD_EN IN_63 NET0279 NAND2_2 
XI432 WORD_EN IN_45 NET0715 NAND2_2 
XI256 WORD_EN IN_1 NET0847 NAND2_2 
XI260 WORD_EN IN_2 NET0645 NAND2_2 
XI284 WORD_EN IN_8 NET0826 NAND2_2 
XI264 WORD_EN IN_3 NET0841 NAND2_2 
XI268 WORD_EN IN_4 NET0633 NAND2_2 
XI288 WORD_EN IN_9 NET0603 NAND2_2 
XI272 WORD_EN IN_5 NET0627 NAND2_2 
XI276 WORD_EN IN_6 NET0621 NAND2_2 
XI296 WORD_EN IN_11 NET0817 NAND2_2 
XI436 WORD_EN IN_46 NET0712 NAND2_2 
XI280 WORD_EN IN_7 NET0829 NAND2_2 
XI308 WORD_EN IN_14 NET0573 NAND2_2 
XI440 WORD_EN IN_47 NET0709 NAND2_2 
XI444 WORD_EN IN_48 NET0369 NAND2_2 
XI312 WORD_EN IN_15 NET0805 NAND2_2 
XI292 WORD_EN IN_10 NET0597 NAND2_2 
XI300 WORD_EN IN_12 NET0585 NAND2_2 
XI304 WORD_EN IN_13 NET0579 NAND2_2 
XI372 WORD_EN IN_30 NET0760 NAND2_2 
XI316 WORD_EN IN_16 NET0561 NAND2_2 
XI376 WORD_EN IN_31 NET0757 NAND2_2 
XI320 WORD_EN IN_17 NET0555 NAND2_2 
XI380 WORD_EN IN_32 NET0754 NAND2_2 
XI324 WORD_EN IN_18 NET0549 NAND2_2 
XI384 WORD_EN IN_33 NET0459 NAND2_2 
XI328 WORD_EN IN_19 NET0543 NAND2_2 
XI388 WORD_EN IN_34 NET0453 NAND2_2 
XI332 WORD_EN IN_20 NET0537 NAND2_2 
XI392 WORD_EN IN_35 NET0745 NAND2_2 
XI336 WORD_EN IN_21 NET0531 NAND2_2 
XI396 WORD_EN IN_36 NET0742 NAND2_2 
XI340 WORD_EN IN_22 NET0525 NAND2_2 
XI400 WORD_EN IN_37 NET0435 NAND2_2 
XI344 WORD_EN IN_23 NET0519 NAND2_2 
XI404 WORD_EN IN_38 NET0429 NAND2_2 
XI348 WORD_EN IN_24 NET0778 NAND2_2 
XI408 WORD_EN IN_39 NET0733 NAND2_2 
XI352 WORD_EN IN_25 NET0775 NAND2_2 
XI412 WORD_EN IN_40 NET0417 NAND2_2 
XI356 WORD_EN IN_26 NET0501 NAND2_2 
XI416 WORD_EN IN_41 NET0727 NAND2_2 
XI360 WORD_EN IN_27 NET0495 NAND2_2 
XI364 WORD_EN IN_28 NET0766 NAND2_2 
XI420 WORD_EN IN_42 NET0405 NAND2_2 
XI424 WORD_EN IN_43 NET0399 NAND2_2 
XI368 WORD_EN IN_29 NET0763 NAND2_2 
XI428 WORD_EN IN_44 NET0718 NAND2_2 
XI0 WORD_EN IN_0 NET50 NAND2_2 
   
   
* FILE NAME: SRAM2_NAND2_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: NAND2.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   OUT = OUT
.SUBCKT NAND2_2 A B OUT 
M3 OUT B VDD! VDD!  PFET  L=200E-9 W=(12.5E-6) AD=+6.25000000E-12 
+AS=+6.25000000E-12 PD=+2.60000000E-05 PS=+2.60000000E-05 NRD=+4.00000000E-02 
+NRS=+4.00000000E-02 M=1.0 
M2 OUT A VDD! VDD!  PFET  L=200E-9 W=(12.5E-6) AD=+6.25000000E-12 
+AS=+6.25000000E-12 PD=+2.60000000E-05 PS=+2.60000000E-05 NRD=+4.00000000E-02 
+NRS=+4.00000000E-02 M=1.0 
M1 OUT A NET15 0  NFET  L=200E-9 W=(8.3E-6) AD=+4.15000000E-12 
+AS=+4.15000000E-12 PD=+1.76000000E-05 PS=+1.76000000E-05 NRD=+6.02409639E-02 
+NRS=+6.02409639E-02 M=1.0 
M0 NET15 B 0 0  NFET  L=200E-9 W=(8.3E-6) AD=+4.15000000E-12 
+AS=+4.15000000E-12 PD=+1.76000000E-05 PS=+1.76000000E-05 NRD=+6.02409639E-02 
+NRS=+6.02409639E-02 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NAND2_2 
* FILE NAME: SRAM2_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_1 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(47.1E-6) AD=+2.35500000E-11 
+AS=+2.35500000E-11 PD=+9.52000000E-05 PS=+9.52000000E-05 NRD=+1.06157113E-02 
+NRS=+1.06157113E-02 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(15.7E-6) AD=+7.85000000E-12 
+AS=+7.85000000E-12 PD=+3.24000000E-05 PS=+3.24000000E-05 NRD=+3.18471338E-02 
+NRS=+3.18471338E-02 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS CONTROL_G19 
* FILE NAME: SRAM2_DUM_SRAM_CELL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: DUM_SRAM_CELL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: BIT = BIT
*                   BIT_STORED = BIT_STORED
*                   WL = WL
*                   BIT_BAR = BIT_BAR
.SUBCKT DUM_SRAM_CELL_G2 BIT BIT_STORED WL BIT_BAR 
M2 BIT_BAR WL VDD! 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M0 BIT_STORED WL BIT 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
XI3 VDD! BIT_STORED INV_1 
XI0 BIT_STORED VDD! INV_1 
   
   
* FILE NAME: SRAM_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_1 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(400E-9) AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(400E-9) AD=+2.00000000E-13 AS=+2.00000000E-13 
+PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 NRS=+1.25000000E+00 
+M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS DUM_SRAM_CELL_G2 
* FILE NAME: SRAM2_PATH1INVS_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: PATH1INVS.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:36 2007.
   
* TERMINAL MAPPING: A_BAR_IN = A_BAR_IN
*                   A_BAR_OUT = A_BAR_OUT
*                   A_IN = A_IN
*                   A_OUT = A_OUT
.SUBCKT PATH1INVS_G5 A_BAR_IN A_BAR_OUT A_IN A_OUT 
XI10 NET014 NET015 INV_1 
XI11 NET015 NET010 INV_2 
XI13 NET010 A_OUT INV_2 
XI6 NET9 NET019 INV_1 
XI4 A_BAR_IN NET9 INV_3 
XI9 NET019 A_BAR_OUT INV_2 
XI0 A_IN NET014 INV_3 
   
   
* FILE NAME: SRAM_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_1 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(32.1E-6) AD=+1.60500000E-11 
+AS=+1.60500000E-11 PD=+6.52000000E-05 PS=+6.52000000E-05 NRD=+1.55763240E-02 
+NRS=+1.55763240E-02 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(10.7E-6) AD=+5.35000000E-12 
+AS=+5.35000000E-12 PD=+2.24000000E-05 PS=+2.24000000E-05 NRD=+4.67289720E-02 
+NRS=+4.67289720E-02 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
* FILE NAME: SRAM_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_3 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(8.5E-6) AD=+4.25000000E-12 
+AS=+4.25000000E-12 PD=+1.80000000E-05 PS=+1.80000000E-05 NRD=+5.88235294E-02 
+NRS=+5.88235294E-02 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(2.8E-6) AD=+1.40000000E-12 AS=+1.40000000E-12 
+PD=+6.60000000E-06 PS=+6.60000000E-06 NRD=+1.78571429E-01 NRS=+1.78571429E-01 
+M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_3 
* FILE NAME: SRAM_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_2 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(121.4E-6) AD=+6.07000000E-11 
+AS=+6.07000000E-11 PD=+2.43800000E-04 PS=+2.43800000E-04 NRD=+4.11861614E-03 
+NRS=+4.11861614E-03 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(40.5E-6) AD=+2.02500000E-11 
+AS=+2.02500000E-11 PD=+8.20000000E-05 PS=+8.20000000E-05 NRD=+1.23456790E-02 
+NRS=+1.23456790E-02 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_2 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS PATH1INVS_G5 
* FILE NAME: SRAM2_TL_PI_MODEL7_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL7.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN<0> = IN_0
*                   IN<1> = IN_1
*                   IN<2> = IN_2
*                   IN<3> = IN_3
*                   IN<4> = IN_4
*                   IN<5> = IN_5
*                   IN<6> = IN_6
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
*                   OUT<3> = OUT_3
*                   OUT<4> = OUT_4
*                   OUT<5> = OUT_5
*                   OUT<6> = OUT_6
.SUBCKT TL_PI_MODEL7_G13 IN_0 IN_1 IN_2 IN_3 IN_4 IN_5 IN_6 OUT_0 OUT_1 OUT_2 
+OUT_3 OUT_4 OUT_5 OUT_6 
XI6 IN_6 OUT_6 TL_PI_MODEL_1 
XI5 IN_5 OUT_5 TL_PI_MODEL_1 
XI4 IN_4 OUT_4 TL_PI_MODEL_1 
XI3 IN_3 OUT_3 TL_PI_MODEL_1 
XI2 IN_2 OUT_2 TL_PI_MODEL_1 
XI1 IN_1 OUT_1 TL_PI_MODEL_1 
XI0 IN_0 OUT_0 TL_PI_MODEL_1 
   
   
* FILE NAME: SRAM2_TL_PI_MODEL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:31 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT TL_PI_MODEL_1 IN OUT 
C0 IN 0  (34E-15) M=1.0 
C1 OUT 0  (34E-15) M=1.0 
R0 IN OUT  (192.0) M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL7_G13 
* FILE NAME: SRAM2_PATH1INVS7_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: PATH1INVS7.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:36 2007.
   
* TERMINAL MAPPING: IN<0> = IN_0
*                   IN<1> = IN_1
*                   IN<2> = IN_2
*                   IN<3> = IN_3
*                   IN<4> = IN_4
*                   IN<5> = IN_5
*                   IN<6> = IN_6
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
*                   OUT<3> = OUT_3
*                   OUT<4> = OUT_4
*                   OUT<5> = OUT_5
*                   OUT<6> = OUT_6
*                   OUT_B<0> = OUT_B_0
*                   OUT_B<1> = OUT_B_1
*                   OUT_B<2> = OUT_B_2
*                   OUT_B<3> = OUT_B_3
*                   OUT_B<4> = OUT_B_4
*                   OUT_B<5> = OUT_B_5
*                   OUT_B<6> = OUT_B_6
.SUBCKT PATH1INVS7_G20 IN_0 IN_1 IN_2 IN_3 IN_4 IN_5 IN_6 OUT_0 OUT_1 OUT_2 
+OUT_3 OUT_4 OUT_5 OUT_6 OUT_B_0 OUT_B_1 OUT_B_2 OUT_B_3 OUT_B_4 OUT_B_5 
+OUT_B_6 
XI6 IN_6 OUT_B_6 IN_6 OUT_6 PATH1INVS_G5 
XI5 IN_5 OUT_B_5 IN_5 OUT_5 PATH1INVS_G5 
XI4 IN_4 OUT_B_4 IN_4 OUT_4 PATH1INVS_G5 
XI3 IN_3 OUT_B_3 IN_3 OUT_3 PATH1INVS_G5 
XI2 IN_2 OUT_B_2 IN_2 OUT_2 PATH1INVS_G5 
XI1 IN_1 OUT_B_1 IN_1 OUT_1 PATH1INVS_G5 
XI0 IN_0 OUT_B_0 IN_0 OUT_0 PATH1INVS_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS PATH1INVS7_G20 
* FILE NAME: SRAM2_COL_DEC_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: COL_DEC.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:35 2007.
   
* TERMINAL MAPPING: ADDRESS<7> = ADDRESS_7
*                   ADDRESS<8> = ADDRESS_8
*                   ADDRESS<9> = ADDRESS_9
*                   ADDRESS_BAR<7> = ADDRESS_BAR_7
*                   ADDRESS_BAR<8> = ADDRESS_BAR_8
*                   ADDRESS_BAR<9> = ADDRESS_BAR_9
*                   ROWDECO<0> = ROWDECO_0
*                   ROWDECO<1> = ROWDECO_1
*                   ROWDECO<2> = ROWDECO_2
*                   ROWDECO<3> = ROWDECO_3
*                   ROWDECO<4> = ROWDECO_4
*                   ROWDECO<5> = ROWDECO_5
*                   ROWDECO<6> = ROWDECO_6
*                   ROWDECO<7> = ROWDECO_7
.SUBCKT COL_DEC_G18 ADDRESS_7 ADDRESS_8 ADDRESS_9 ADDRESS_BAR_7 ADDRESS_BAR_8 
+ADDRESS_BAR_9 ROWDECO_0 ROWDECO_1 ROWDECO_2 ROWDECO_3 ROWDECO_4 ROWDECO_5 
+ROWDECO_6 ROWDECO_7 
XI0 ROWDECO_0 ROWDECO_1 ROWDECO_2 ROWDECO_3 ROWDECO_4 ROWDECO_5 ROWDECO_6 
+ROWDECO_7 ADDRESS_7 ADDRESS_8 ADDRESS_9 ADDRESS_BAR_7 ADDRESS_BAR_8 
+ADDRESS_BAR_9 VDD! RDEC3TO8A_G4 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS COL_DEC_G18 
* FILE NAME: SRAM2_REG32_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: REG32.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:42 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   IN<0> = IN_0
*                   IN<1> = IN_1
*                   IN<2> = IN_2
*                   IN<3> = IN_3
*                   IN<4> = IN_4
*                   IN<5> = IN_5
*                   IN<6> = IN_6
*                   IN<7> = IN_7
*                   IN<8> = IN_8
*                   IN<9> = IN_9
*                   IN<10> = IN_10
*                   IN<11> = IN_11
*                   IN<12> = IN_12
*                   IN<13> = IN_13
*                   IN<14> = IN_14
*                   IN<15> = IN_15
*                   IN<16> = IN_16
*                   IN<17> = IN_17
*                   IN<18> = IN_18
*                   IN<19> = IN_19
*                   IN<20> = IN_20
*                   IN<21> = IN_21
*                   IN<22> = IN_22
*                   IN<23> = IN_23
*                   IN<24> = IN_24
*                   IN<25> = IN_25
*                   IN<26> = IN_26
*                   IN<27> = IN_27
*                   IN<28> = IN_28
*                   IN<29> = IN_29
*                   IN<30> = IN_30
*                   IN<31> = IN_31
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
*                   OUT<3> = OUT_3
*                   OUT<4> = OUT_4
*                   OUT<5> = OUT_5
*                   OUT<6> = OUT_6
*                   OUT<7> = OUT_7
*                   OUT<8> = OUT_8
*                   OUT<9> = OUT_9
*                   OUT<10> = OUT_10
*                   OUT<11> = OUT_11
*                   OUT<12> = OUT_12
*                   OUT<13> = OUT_13
*                   OUT<14> = OUT_14
*                   OUT<15> = OUT_15
*                   OUT<16> = OUT_16
*                   OUT<17> = OUT_17
*                   OUT<18> = OUT_18
*                   OUT<19> = OUT_19
*                   OUT<20> = OUT_20
*                   OUT<21> = OUT_21
*                   OUT<22> = OUT_22
*                   OUT<23> = OUT_23
*                   OUT<24> = OUT_24
*                   OUT<25> = OUT_25
*                   OUT<26> = OUT_26
*                   OUT<27> = OUT_27
*                   OUT<28> = OUT_28
*                   OUT<29> = OUT_29
*                   OUT<30> = OUT_30
*                   OUT<31> = OUT_31
.SUBCKT REG32_G24 CLK IN_0 IN_1 IN_2 IN_3 IN_4 IN_5 IN_6 IN_7 IN_8 IN_9 IN_10 
+IN_11 IN_12 IN_13 IN_14 IN_15 IN_16 IN_17 IN_18 IN_19 IN_20 IN_21 IN_22 IN_23 
+IN_24 IN_25 IN_26 IN_27 IN_28 IN_29 IN_30 IN_31 OUT_0 OUT_1 OUT_2 OUT_3 OUT_4 
+OUT_5 OUT_6 OUT_7 OUT_8 OUT_9 OUT_10 OUT_11 OUT_12 OUT_13 OUT_14 OUT_15 OUT_16 
+OUT_17 OUT_18 OUT_19 OUT_20 OUT_21 OUT_22 OUT_23 OUT_24 OUT_25 OUT_26 OUT_27 
+OUT_28 OUT_29 OUT_30 OUT_31 
XI31 CLK IN_31 OUT_31 DFFPOSX1_G6 
XI30 CLK IN_30 OUT_30 DFFPOSX1_G6 
XI29 CLK IN_29 OUT_29 DFFPOSX1_G6 
XI28 CLK IN_28 OUT_28 DFFPOSX1_G6 
XI27 CLK IN_27 OUT_27 DFFPOSX1_G6 
XI26 CLK IN_26 OUT_26 DFFPOSX1_G6 
XI25 CLK IN_25 OUT_25 DFFPOSX1_G6 
XI24 CLK IN_24 OUT_24 DFFPOSX1_G6 
XI23 CLK IN_23 OUT_23 DFFPOSX1_G6 
XI22 CLK IN_22 OUT_22 DFFPOSX1_G6 
XI21 CLK IN_21 OUT_21 DFFPOSX1_G6 
XI20 CLK IN_20 OUT_20 DFFPOSX1_G6 
XI19 CLK IN_19 OUT_19 DFFPOSX1_G6 
XI18 CLK IN_18 OUT_18 DFFPOSX1_G6 
XI17 CLK IN_17 OUT_17 DFFPOSX1_G6 
XI16 CLK IN_16 OUT_16 DFFPOSX1_G6 
XI15 CLK IN_15 OUT_15 DFFPOSX1_G6 
XI14 CLK IN_14 OUT_14 DFFPOSX1_G6 
XI13 CLK IN_13 OUT_13 DFFPOSX1_G6 
XI12 CLK IN_12 OUT_12 DFFPOSX1_G6 
XI11 CLK IN_11 OUT_11 DFFPOSX1_G6 
XI10 CLK IN_10 OUT_10 DFFPOSX1_G6 
XI9 CLK IN_9 OUT_9 DFFPOSX1_G6 
XI8 CLK IN_8 OUT_8 DFFPOSX1_G6 
XI7 CLK IN_7 OUT_7 DFFPOSX1_G6 
XI6 CLK IN_6 OUT_6 DFFPOSX1_G6 
XI5 CLK IN_5 OUT_5 DFFPOSX1_G6 
XI4 CLK IN_4 OUT_4 DFFPOSX1_G6 
XI3 CLK IN_3 OUT_3 DFFPOSX1_G6 
XI2 CLK IN_2 OUT_2 DFFPOSX1_G6 
XI1 CLK IN_1 OUT_1 DFFPOSX1_G6 
XI0 CLK IN_0 OUT_0 DFFPOSX1_G6 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS REG32_G24 
* FILE NAME: SRAM2_SRAM_CELL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SRAM_CELL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: BIT = BIT
*                   BIT_BAR_STORED = BIT_BAR_STORED
*                   BIT_STORED = BIT_STORED
*                   WL = WL
*                   BIT_BAR = BIT_BAR
.SUBCKT SRAM_CELL_G1 BIT BIT_BAR_STORED BIT_STORED WL BIT_BAR 
M2 BIT_BAR WL BIT_BAR_STORED 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M0 BIT_STORED WL BIT 0  NFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
XI3 BIT_BAR_STORED BIT_STORED INV_1 
XI0 BIT_STORED BIT_BAR_STORED INV_1 
   
   
* FILE NAME: SRAM_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_1 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(400E-9) AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(400E-9) AD=+2.00000000E-13 AS=+2.00000000E-13 
+PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 NRS=+1.25000000E+00 
+M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SRAM_CELL_G1 
* FILE NAME: OSU_STDCELLS_DFFPOSX1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: DFFPOSX1.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D = D
*                   Q = Q
.SUBCKT DFFPOSX1_G6 CLK D Q 
M64 NET071 NET33 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M58 NET33 CLK NET18 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M57 CLK_B CLK 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M61 NET18 NET071 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M60 Q NET27 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M66 NET24 NET071 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M65 NET27 CLK NET24 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M67 NET9 Q 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 PS=3E-6 
+M=1 
M62 NET33 CLK_B NET30 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 
+PD=3E-6 PS=3E-6 M=1 
M59 NET27 CLK_B NET9 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M63 NET30 D 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M46 CLK_B CLK VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M47 NET50 NET071 VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M48 NET41 Q VDD! VDD!  TSMC20P  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M49 Q NET27 VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M50 NET33 CLK_B NET50 VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M51 NET62 D VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M52 NET33 CLK NET62 VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M53 NET56 NET071 VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M54 NET27 CLK_B NET56 VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M55 NET071 NET33 VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M56 NET27 CLK NET41 VDD!  TSMC20P  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 
+PD=3E-6 PS=3E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS DFFPOSX1_G6 
* FILE NAME: SRAM2_RDEC7TO128_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: RDEC7TO128.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:39 2007.
   
* TERMINAL MAPPING: RDECO<0> = RDECO_0
*                   RDECO<1> = RDECO_1
*                   RDECO<2> = RDECO_2
*                   RDECO<3> = RDECO_3
*                   RDECO<4> = RDECO_4
*                   RDECO<5> = RDECO_5
*                   RDECO<6> = RDECO_6
*                   RDECO<7> = RDECO_7
*                   RDECO<8> = RDECO_8
*                   RDECO<9> = RDECO_9
*                   RDECO<10> = RDECO_10
*                   RDECO<11> = RDECO_11
*                   RDECO<12> = RDECO_12
*                   RDECO<13> = RDECO_13
*                   RDECO<14> = RDECO_14
*                   RDECO<15> = RDECO_15
*                   RDECO<16> = RDECO_16
*                   RDECO<17> = RDECO_17
*                   RDECO<18> = RDECO_18
*                   RDECO<19> = RDECO_19
*                   RDECO<20> = RDECO_20
*                   RDECO<21> = RDECO_21
*                   RDECO<22> = RDECO_22
*                   RDECO<23> = RDECO_23
*                   RDECO<24> = RDECO_24
*                   RDECO<25> = RDECO_25
*                   RDECO<26> = RDECO_26
*                   RDECO<27> = RDECO_27
*                   RDECO<28> = RDECO_28
*                   RDECO<29> = RDECO_29
*                   RDECO<30> = RDECO_30
*                   RDECO<31> = RDECO_31
*                   RDECO<32> = RDECO_32
*                   RDECO<33> = RDECO_33
*                   RDECO<34> = RDECO_34
*                   RDECO<35> = RDECO_35
*                   RDECO<36> = RDECO_36
*                   RDECO<37> = RDECO_37
*                   RDECO<38> = RDECO_38
*                   RDECO<39> = RDECO_39
*                   RDECO<40> = RDECO_40
*                   RDECO<41> = RDECO_41
*                   RDECO<42> = RDECO_42
*                   RDECO<43> = RDECO_43
*                   RDECO<44> = RDECO_44
*                   RDECO<45> = RDECO_45
*                   RDECO<46> = RDECO_46
*                   RDECO<47> = RDECO_47
*                   RDECO<48> = RDECO_48
*                   RDECO<49> = RDECO_49
*                   RDECO<50> = RDECO_50
*                   RDECO<51> = RDECO_51
*                   RDECO<52> = RDECO_52
*                   RDECO<53> = RDECO_53
*                   RDECO<54> = RDECO_54
*                   RDECO<55> = RDECO_55
*                   RDECO<56> = RDECO_56
*                   RDECO<57> = RDECO_57
*                   RDECO<58> = RDECO_58
*                   RDECO<59> = RDECO_59
*                   RDECO<60> = RDECO_60
*                   RDECO<61> = RDECO_61
*                   RDECO<62> = RDECO_62
*                   RDECO<63> = RDECO_63
*                   RDECO<64> = RDECO_64
*                   RDECO<65> = RDECO_65
*                   RDECO<66> = RDECO_66
*                   RDECO<67> = RDECO_67
*                   RDECO<68> = RDECO_68
*                   RDECO<69> = RDECO_69
*                   RDECO<70> = RDECO_70
*                   RDECO<71> = RDECO_71
*                   RDECO<72> = RDECO_72
*                   RDECO<73> = RDECO_73
*                   RDECO<74> = RDECO_74
*                   RDECO<75> = RDECO_75
*                   RDECO<76> = RDECO_76
*                   RDECO<77> = RDECO_77
*                   RDECO<78> = RDECO_78
*                   RDECO<79> = RDECO_79
*                   RDECO<80> = RDECO_80
*                   RDECO<81> = RDECO_81
*                   RDECO<82> = RDECO_82
*                   RDECO<83> = RDECO_83
*                   RDECO<84> = RDECO_84
*                   RDECO<85> = RDECO_85
*                   RDECO<86> = RDECO_86
*                   RDECO<87> = RDECO_87
*                   RDECO<88> = RDECO_88
*                   RDECO<89> = RDECO_89
*                   RDECO<90> = RDECO_90
*                   RDECO<91> = RDECO_91
*                   RDECO<92> = RDECO_92
*                   RDECO<93> = RDECO_93
*                   RDECO<94> = RDECO_94
*                   RDECO<95> = RDECO_95
*                   RDECO<96> = RDECO_96
*                   RDECO<97> = RDECO_97
*                   RDECO<98> = RDECO_98
*                   RDECO<99> = RDECO_99
*                   RDECO<100> = RDECO_100
*                   RDECO<101> = RDECO_101
*                   RDECO<102> = RDECO_102
*                   RDECO<103> = RDECO_103
*                   RDECO<104> = RDECO_104
*                   RDECO<105> = RDECO_105
*                   RDECO<106> = RDECO_106
*                   RDECO<107> = RDECO_107
*                   RDECO<108> = RDECO_108
*                   RDECO<109> = RDECO_109
*                   RDECO<110> = RDECO_110
*                   RDECO<111> = RDECO_111
*                   RDECO<112> = RDECO_112
*                   RDECO<113> = RDECO_113
*                   RDECO<114> = RDECO_114
*                   RDECO<115> = RDECO_115
*                   RDECO<116> = RDECO_116
*                   RDECO<117> = RDECO_117
*                   RDECO<118> = RDECO_118
*                   RDECO<119> = RDECO_119
*                   RDECO<120> = RDECO_120
*                   RDECO<121> = RDECO_121
*                   RDECO<122> = RDECO_122
*                   RDECO<123> = RDECO_123
*                   RDECO<124> = RDECO_124
*                   RDECO<125> = RDECO_125
*                   RDECO<126> = RDECO_126
*                   RDECO<127> = RDECO_127
*                   RI<0> = RI_0
*                   RI<1> = RI_1
*                   RI<2> = RI_2
*                   RI<3> = RI_3
*                   RI<4> = RI_4
*                   RI<5> = RI_5
*                   RI<6> = RI_6
*                   RIB<0> = RIB_0
*                   RIB<1> = RIB_1
*                   RIB<2> = RIB_2
*                   RIB<3> = RIB_3
*                   RIB<4> = RIB_4
*                   RIB<5> = RIB_5
*                   RIB<6> = RIB_6
.SUBCKT RDEC7TO128_G22 RDECO_0 RDECO_1 RDECO_2 RDECO_3 RDECO_4 RDECO_5 RDECO_6 
+RDECO_7 RDECO_8 RDECO_9 RDECO_10 RDECO_11 RDECO_12 RDECO_13 RDECO_14 RDECO_15 
+RDECO_16 RDECO_17 RDECO_18 RDECO_19 RDECO_20 RDECO_21 RDECO_22 RDECO_23 
+RDECO_24 RDECO_25 RDECO_26 RDECO_27 RDECO_28 RDECO_29 RDECO_30 RDECO_31 
+RDECO_32 RDECO_33 RDECO_34 RDECO_35 RDECO_36 RDECO_37 RDECO_38 RDECO_39 
+RDECO_40 RDECO_41 RDECO_42 RDECO_43 RDECO_44 RDECO_45 RDECO_46 RDECO_47 
+RDECO_48 RDECO_49 RDECO_50 RDECO_51 RDECO_52 RDECO_53 RDECO_54 RDECO_55 
+RDECO_56 RDECO_57 RDECO_58 RDECO_59 RDECO_60 RDECO_61 RDECO_62 RDECO_63 
+RDECO_64 RDECO_65 RDECO_66 RDECO_67 RDECO_68 RDECO_69 RDECO_70 RDECO_71 
+RDECO_72 RDECO_73 RDECO_74 RDECO_75 RDECO_76 RDECO_77 RDECO_78 RDECO_79 
+RDECO_80 RDECO_81 RDECO_82 RDECO_83 RDECO_84 RDECO_85 RDECO_86 RDECO_87 
+RDECO_88 RDECO_89 RDECO_90 RDECO_91 RDECO_92 RDECO_93 RDECO_94 RDECO_95 
+RDECO_96 RDECO_97 RDECO_98 RDECO_99 RDECO_100 RDECO_101 RDECO_102 RDECO_103 
+RDECO_104 RDECO_105 RDECO_106 RDECO_107 RDECO_108 RDECO_109 RDECO_110 
+RDECO_111 RDECO_112 RDECO_113 RDECO_114 RDECO_115 RDECO_116 RDECO_117 
+RDECO_118 RDECO_119 RDECO_120 RDECO_121 RDECO_122 RDECO_123 RDECO_124 
+RDECO_125 RDECO_126 RDECO_127 RI_0 RI_1 RI_2 RI_3 RI_4 RI_5 RI_6 RIB_0 RIB_1 
+RIB_2 RIB_3 RIB_4 RIB_5 RIB_6 
M128 RDECO_64 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M127 RDECO_65 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M126 RDECO_66 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M125 RDECO_67 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M124 RDECO_68 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M123 RDECO_69 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M122 RDECO_70 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M121 RDECO_71 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M120 RDECO_72 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M119 RDECO_73 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M118 RDECO_74 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M117 RDECO_75 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M116 RDECO_76 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M115 RDECO_77 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M114 RDECO_78 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M113 RDECO_79 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M112 RDECO_80 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M111 RDECO_81 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M110 RDECO_82 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M109 RDECO_83 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M108 RDECO_84 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M107 RDECO_85 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M106 RDECO_86 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M105 RDECO_87 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M104 RDECO_88 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M103 RDECO_89 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M102 RDECO_90 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M101 RDECO_91 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M100 RDECO_92 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M99 RDECO_93 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M98 RDECO_94 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M97 RDECO_95 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M96 RDECO_96 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M95 RDECO_97 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M94 RDECO_98 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M93 RDECO_99 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M92 RDECO_100 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M91 RDECO_101 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M90 RDECO_102 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M89 RDECO_103 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M88 RDECO_104 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M87 RDECO_105 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M86 RDECO_106 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M85 RDECO_107 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M84 RDECO_108 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M83 RDECO_109 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M82 RDECO_110 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M81 RDECO_111 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M80 RDECO_112 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M79 RDECO_113 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M78 RDECO_114 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M77 RDECO_115 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M76 RDECO_116 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M75 RDECO_117 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M74 RDECO_118 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M73 RDECO_119 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M72 RDECO_120 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M71 RDECO_121 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M70 RDECO_122 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M69 RDECO_123 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M68 RDECO_124 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M67 RDECO_125 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M66 RDECO_126 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M65 RDECO_127 RIB_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M64 RDECO_63 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M63 RDECO_62 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M62 RDECO_61 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M61 RDECO_60 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M60 RDECO_59 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M59 RDECO_58 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M58 RDECO_57 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M57 RDECO_56 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M56 RDECO_55 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M55 RDECO_54 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M54 RDECO_53 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M53 RDECO_52 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M52 RDECO_51 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M51 RDECO_50 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M50 RDECO_49 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M49 RDECO_48 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M48 RDECO_47 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M47 RDECO_46 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M46 RDECO_45 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M45 RDECO_44 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M44 RDECO_43 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M43 RDECO_42 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M42 RDECO_41 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M41 RDECO_40 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M40 RDECO_39 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M39 RDECO_38 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M38 RDECO_37 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M37 RDECO_36 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M36 RDECO_35 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M35 RDECO_34 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M34 RDECO_33 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M33 RDECO_32 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M30 RDECO_29 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M29 RDECO_28 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M28 RDECO_27 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M27 RDECO_26 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M26 RDECO_25 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M25 RDECO_24 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M24 RDECO_23 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M23 RDECO_22 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M22 RDECO_21 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M21 RDECO_20 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M20 RDECO_19 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M19 RDECO_18 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M18 RDECO_17 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M17 RDECO_16 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M16 RDECO_15 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M15 RDECO_14 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M14 RDECO_13 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M13 RDECO_12 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M12 RDECO_11 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M11 RDECO_10 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M10 RDECO_9 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M9 RDECO_8 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M8 RDECO_7 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M7 RDECO_6 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M6 RDECO_5 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M5 RDECO_4 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M4 RDECO_3 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M3 RDECO_2 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M2 RDECO_1 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M1 RDECO_0 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M31 RDECO_30 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M32 RDECO_31 RI_6 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M129 NET4 RIB_6 VDD! VDD!  PFET  L=200E-9 W=294.4E-6 AD=+1.47200000E-10 
+AS=+1.47200000E-10 PD=+5.89800000E-04 PS=+5.89800000E-04 NRD=+1.69836957E-03 
+NRS=+1.69836957E-03 M=1.0 
M0 NET81 RI_6 VDD! VDD!  PFET  L=200E-9 W=294.4E-6 AD=+1.47200000E-10 
+AS=+1.47200000E-10 PD=+5.89800000E-04 PS=+5.89800000E-04 NRD=+1.69836957E-03 
+NRS=+1.69836957E-03 M=1.0 
XI1 RDECO_64 RDECO_65 RDECO_66 RDECO_67 RDECO_68 RDECO_69 RDECO_70 RDECO_71 
+RDECO_72 RDECO_73 RDECO_74 RDECO_75 RDECO_76 RDECO_77 RDECO_78 RDECO_79 
+RDECO_80 RDECO_81 RDECO_82 RDECO_83 RDECO_84 RDECO_85 RDECO_86 RDECO_87 
+RDECO_88 RDECO_89 RDECO_90 RDECO_91 RDECO_92 RDECO_93 RDECO_94 RDECO_95 
+RDECO_96 RDECO_97 RDECO_98 RDECO_99 RDECO_100 RDECO_101 RDECO_102 RDECO_103 
+RDECO_104 RDECO_105 RDECO_106 RDECO_107 RDECO_108 RDECO_109 RDECO_110 
+RDECO_111 RDECO_112 RDECO_113 RDECO_114 RDECO_115 RDECO_116 RDECO_117 
+RDECO_118 RDECO_119 RDECO_120 RDECO_121 RDECO_122 RDECO_123 RDECO_124 
+RDECO_125 RDECO_126 RDECO_127 RI_0 RI_1 RI_2 RI_3 RI_4 RI_5 RIB_0 RIB_1 RIB_2 
+RIB_3 RIB_4 RIB_5 NET4 RDEC6TO64_G10 
XI0 RDECO_0 RDECO_1 RDECO_2 RDECO_3 RDECO_4 RDECO_5 RDECO_6 RDECO_7 RDECO_8 
+RDECO_9 RDECO_10 RDECO_11 RDECO_12 RDECO_13 RDECO_14 RDECO_15 RDECO_16 
+RDECO_17 RDECO_18 RDECO_19 RDECO_20 RDECO_21 RDECO_22 RDECO_23 RDECO_24 
+RDECO_25 RDECO_26 RDECO_27 RDECO_28 RDECO_29 RDECO_30 RDECO_31 RDECO_32 
+RDECO_33 RDECO_34 RDECO_35 RDECO_36 RDECO_37 RDECO_38 RDECO_39 RDECO_40 
+RDECO_41 RDECO_42 RDECO_43 RDECO_44 RDECO_45 RDECO_46 RDECO_47 RDECO_48 
+RDECO_49 RDECO_50 RDECO_51 RDECO_52 RDECO_53 RDECO_54 RDECO_55 RDECO_56 
+RDECO_57 RDECO_58 RDECO_59 RDECO_60 RDECO_61 RDECO_62 RDECO_63 RI_0 RI_1 RI_2 
+RI_3 RI_4 RI_5 RIB_0 RIB_1 RIB_2 RIB_3 RIB_4 RIB_5 NET81 RDEC6TO64_G10 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS RDEC7TO128_G22 
* FILE NAME: SRAM_RDEC5TO32_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: RDEC5TO32.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:38 2007.
   
* TERMINAL MAPPING: RDECO<0> = RDECO_0
*                   RDECO<1> = RDECO_1
*                   RDECO<2> = RDECO_2
*                   RDECO<3> = RDECO_3
*                   RDECO<4> = RDECO_4
*                   RDECO<5> = RDECO_5
*                   RDECO<6> = RDECO_6
*                   RDECO<7> = RDECO_7
*                   RDECO<8> = RDECO_8
*                   RDECO<9> = RDECO_9
*                   RDECO<10> = RDECO_10
*                   RDECO<11> = RDECO_11
*                   RDECO<12> = RDECO_12
*                   RDECO<13> = RDECO_13
*                   RDECO<14> = RDECO_14
*                   RDECO<15> = RDECO_15
*                   RDECO<16> = RDECO_16
*                   RDECO<17> = RDECO_17
*                   RDECO<18> = RDECO_18
*                   RDECO<19> = RDECO_19
*                   RDECO<20> = RDECO_20
*                   RDECO<21> = RDECO_21
*                   RDECO<22> = RDECO_22
*                   RDECO<23> = RDECO_23
*                   RDECO<24> = RDECO_24
*                   RDECO<25> = RDECO_25
*                   RDECO<26> = RDECO_26
*                   RDECO<27> = RDECO_27
*                   RDECO<28> = RDECO_28
*                   RDECO<29> = RDECO_29
*                   RDECO<30> = RDECO_30
*                   RDECO<31> = RDECO_31
*                   RI<0> = RI_0
*                   RI<1> = RI_1
*                   RI<2> = RI_2
*                   RI<3> = RI_3
*                   RI<4> = RI_4
*                   RIB<0> = RIB_0
*                   RIB<1> = RIB_1
*                   RIB<2> = RIB_2
*                   RIB<3> = RIB_3
*                   RIB<4> = RIB_4
*                   TOP = TOP
.SUBCKT RDEC5TO32_G9 RDECO_0 RDECO_1 RDECO_2 RDECO_3 RDECO_4 RDECO_5 RDECO_6 
+RDECO_7 RDECO_8 RDECO_9 RDECO_10 RDECO_11 RDECO_12 RDECO_13 RDECO_14 RDECO_15 
+RDECO_16 RDECO_17 RDECO_18 RDECO_19 RDECO_20 RDECO_21 RDECO_22 RDECO_23 
+RDECO_24 RDECO_25 RDECO_26 RDECO_27 RDECO_28 RDECO_29 RDECO_30 RDECO_31 RI_0 
+RI_1 RI_2 RI_3 RI_4 RIB_0 RIB_1 RIB_2 RIB_3 RIB_4 TOP 
XI3 RDECO_0 RDECO_1 RDECO_2 RDECO_3 RDECO_4 RDECO_5 RDECO_6 RDECO_7 RDECO_8 
+RDECO_9 RDECO_10 RDECO_11 RDECO_12 RDECO_13 RDECO_14 RDECO_15 RI_0 RI_1 RI_2 
+RI_3 RIB_0 RIB_1 RIB_2 RIB_3 NET32 RDEC4TO16A_G8 
XI4 RDECO_16 RDECO_17 RDECO_18 RDECO_19 RDECO_20 RDECO_21 RDECO_22 RDECO_23 
+RDECO_24 RDECO_25 RDECO_26 RDECO_27 RDECO_28 RDECO_29 RDECO_30 RDECO_31 RI_0 
+RI_1 RI_2 RI_3 RIB_0 RIB_1 RIB_2 RIB_3 NET7 RDEC4TO16A_G8 
M33 RDECO_31 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M32 RDECO_30 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M31 RDECO_29 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M30 RDECO_28 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M29 RDECO_27 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M28 RDECO_26 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M27 RDECO_25 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M26 RDECO_24 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M25 RDECO_23 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M24 RDECO_22 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M23 RDECO_21 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M22 RDECO_20 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M21 RDECO_19 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M20 RDECO_18 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M19 RDECO_17 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M18 RDECO_16 RIB_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M17 RDECO_15 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M16 RDECO_14 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M15 RDECO_13 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M14 RDECO_12 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M13 RDECO_11 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M12 RDECO_10 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M11 RDECO_9 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M10 RDECO_8 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M9 RDECO_7 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M8 RDECO_6 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M7 RDECO_5 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M6 RDECO_4 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M5 RDECO_3 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M4 RDECO_2 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M3 RDECO_1 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M2 RDECO_0 RI_4 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M1 NET7 RIB_4 TOP VDD!  PFET  L=200E-9 W=73.6E-6 AD=+3.68000000E-11 
+AS=+3.68000000E-11 PD=+1.48200000E-04 PS=+1.48200000E-04 NRD=+6.79347826E-03 
+NRS=+6.79347826E-03 M=1.0 
M0 NET32 RI_4 TOP VDD!  PFET  L=200E-9 W=73.6E-6 AD=+3.68000000E-11 
+AS=+3.68000000E-11 PD=+1.48200000E-04 PS=+1.48200000E-04 NRD=+6.79347826E-03 
+NRS=+6.79347826E-03 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS RDEC5TO32_G9 
* FILE NAME: SRAM2_INV32_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV32.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:41 2007.
   
* TERMINAL MAPPING: IN<0> = IN_0
*                   IN<1> = IN_1
*                   IN<2> = IN_2
*                   IN<3> = IN_3
*                   IN<4> = IN_4
*                   IN<5> = IN_5
*                   IN<6> = IN_6
*                   IN<7> = IN_7
*                   IN<8> = IN_8
*                   IN<9> = IN_9
*                   IN<10> = IN_10
*                   IN<11> = IN_11
*                   IN<12> = IN_12
*                   IN<13> = IN_13
*                   IN<14> = IN_14
*                   IN<15> = IN_15
*                   IN<16> = IN_16
*                   IN<17> = IN_17
*                   IN<18> = IN_18
*                   IN<19> = IN_19
*                   IN<20> = IN_20
*                   IN<21> = IN_21
*                   IN<22> = IN_22
*                   IN<23> = IN_23
*                   IN<24> = IN_24
*                   IN<25> = IN_25
*                   IN<26> = IN_26
*                   IN<27> = IN_27
*                   IN<28> = IN_28
*                   IN<29> = IN_29
*                   IN<30> = IN_30
*                   IN<31> = IN_31
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
*                   OUT<3> = OUT_3
*                   OUT<4> = OUT_4
*                   OUT<5> = OUT_5
*                   OUT<6> = OUT_6
*                   OUT<7> = OUT_7
*                   OUT<8> = OUT_8
*                   OUT<9> = OUT_9
*                   OUT<10> = OUT_10
*                   OUT<11> = OUT_11
*                   OUT<12> = OUT_12
*                   OUT<13> = OUT_13
*                   OUT<14> = OUT_14
*                   OUT<15> = OUT_15
*                   OUT<16> = OUT_16
*                   OUT<17> = OUT_17
*                   OUT<18> = OUT_18
*                   OUT<19> = OUT_19
*                   OUT<20> = OUT_20
*                   OUT<21> = OUT_21
*                   OUT<22> = OUT_22
*                   OUT<23> = OUT_23
*                   OUT<24> = OUT_24
*                   OUT<25> = OUT_25
*                   OUT<26> = OUT_26
*                   OUT<27> = OUT_27
*                   OUT<28> = OUT_28
*                   OUT<29> = OUT_29
*                   OUT<30> = OUT_30
*                   OUT<31> = OUT_31
.SUBCKT INV32_G23 IN_0 IN_1 IN_2 IN_3 IN_4 IN_5 IN_6 IN_7 IN_8 IN_9 IN_10 
+IN_11 IN_12 IN_13 IN_14 IN_15 IN_16 IN_17 IN_18 IN_19 IN_20 IN_21 IN_22 IN_23 
+IN_24 IN_25 IN_26 IN_27 IN_28 IN_29 IN_30 IN_31 OUT_0 OUT_1 OUT_2 OUT_3 OUT_4 
+OUT_5 OUT_6 OUT_7 OUT_8 OUT_9 OUT_10 OUT_11 OUT_12 OUT_13 OUT_14 OUT_15 OUT_16 
+OUT_17 OUT_18 OUT_19 OUT_20 OUT_21 OUT_22 OUT_23 OUT_24 OUT_25 OUT_26 OUT_27 
+OUT_28 OUT_29 OUT_30 OUT_31 
XI31 IN_31 OUT_31 INV_1 
XI30 IN_30 OUT_30 INV_1 
XI29 IN_29 OUT_29 INV_1 
XI28 IN_28 OUT_28 INV_1 
XI27 IN_27 OUT_27 INV_1 
XI26 IN_26 OUT_26 INV_1 
XI25 IN_25 OUT_25 INV_1 
XI24 IN_24 OUT_24 INV_1 
XI23 IN_23 OUT_23 INV_1 
XI22 IN_22 OUT_22 INV_1 
XI21 IN_21 OUT_21 INV_1 
XI20 IN_20 OUT_20 INV_1 
XI19 IN_19 OUT_19 INV_1 
XI18 IN_18 OUT_18 INV_1 
XI17 IN_17 OUT_17 INV_1 
XI16 IN_16 OUT_16 INV_1 
XI15 IN_15 OUT_15 INV_1 
XI14 IN_14 OUT_14 INV_1 
XI13 IN_13 OUT_13 INV_1 
XI12 IN_12 OUT_12 INV_1 
XI11 IN_11 OUT_11 INV_1 
XI10 IN_10 OUT_10 INV_1 
XI9 IN_9 OUT_9 INV_1 
XI8 IN_8 OUT_8 INV_1 
XI7 IN_7 OUT_7 INV_1 
XI6 IN_6 OUT_6 INV_1 
XI5 IN_5 OUT_5 INV_1 
XI4 IN_4 OUT_4 INV_1 
XI3 IN_3 OUT_3 INV_1 
XI2 IN_2 OUT_2 INV_1 
XI1 IN_1 OUT_1 INV_1 
XI0 IN_0 OUT_0 INV_1 
   
   
* FILE NAME: SRAM2_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_1 IN OUT 
M1 OUT IN VDD! VDD!  PFET  L=200E-9 W=(1.2E-6) AD=+6.00000000E-13 
+AS=+6.00000000E-13 PD=+3.40000000E-06 PS=+3.40000000E-06 NRD=+4.16666667E-01 
+NRS=+4.16666667E-01 M=1.0 
M0 OUT IN 0 0  NFET  L=200E-9 W=(400E-9) AD=+2.00000000E-13 AS=+2.00000000E-13 
+PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 NRS=+1.25000000E+00 
+M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV32_G23 
* FILE NAME: SRAM2_TL_PI_MODEL3_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL3.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN<0> = IN_0
*                   IN<1> = IN_1
*                   IN<2> = IN_2
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
.SUBCKT TL_PI_MODEL3_G14 IN_0 IN_1 IN_2 OUT_0 OUT_1 OUT_2 
XI2 IN_2 OUT_2 TL_PI_MODEL_1 
XI1 IN_1 OUT_1 TL_PI_MODEL_1 
XI0 IN_0 OUT_0 TL_PI_MODEL_1 
   
   
* FILE NAME: SRAM2_TL_PI_MODEL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:31 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT TL_PI_MODEL_1 IN OUT 
C0 IN 0  (33E-15) M=1.0 
C1 OUT 0  (33E-15) M=1.0 
R0 IN OUT  (128.0) M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL3_G14 
* FILE NAME: SRAM_RDEC3TO8A_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: RDEC3TO8A.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:37 2007.
   
* TERMINAL MAPPING: RDECO<0> = RDECO_0
*                   RDECO<1> = RDECO_1
*                   RDECO<2> = RDECO_2
*                   RDECO<3> = RDECO_3
*                   RDECO<4> = RDECO_4
*                   RDECO<5> = RDECO_5
*                   RDECO<6> = RDECO_6
*                   RDECO<7> = RDECO_7
*                   RI<0> = RI_0
*                   RI<1> = RI_1
*                   RI<2> = RI_2
*                   RIB<0> = RIB_0
*                   RIB<1> = RIB_1
*                   RIB<2> = RIB_2
*                   TOP = TOP
.SUBCKT RDEC3TO8A_G7 RDECO_0 RDECO_1 RDECO_2 RDECO_3 RDECO_4 RDECO_5 RDECO_6 
+RDECO_7 RI_0 RI_1 RI_2 RIB_0 RIB_1 RIB_2 TOP 
M37 NET0174 RIB_2 TOP VDD!  PFET  L=200E-9 W=16.4E-6 AD=+8.20000000E-12 
+AS=+8.20000000E-12 PD=+3.38000000E-05 PS=+3.38000000E-05 NRD=+3.04878049E-02 
+NRS=+3.04878049E-02 M=1.0 
M36 NET0175 RI_2 TOP VDD!  PFET  L=200E-9 W=16.4E-6 AD=+8.20000000E-12 
+AS=+8.20000000E-12 PD=+3.38000000E-05 PS=+3.38000000E-05 NRD=+3.04878049E-02 
+NRS=+3.04878049E-02 M=1.0 
M28 RDECO_1 RIB_0 NET056 VDD!  PFET  L=200E-9 W=4.1E-6 AD=+2.05000000E-12 
+AS=+2.05000000E-12 PD=+9.20000000E-06 PS=+9.20000000E-06 NRD=+1.21951220E-01 
+NRS=+1.21951220E-01 M=1.0 
M29 RDECO_3 RIB_0 NET068 VDD!  PFET  L=200E-9 W=4.1E-6 AD=+2.05000000E-12 
+AS=+2.05000000E-12 PD=+9.20000000E-06 PS=+9.20000000E-06 NRD=+1.21951220E-01 
+NRS=+1.21951220E-01 M=1.0 
M30 RDECO_5 RIB_0 NET050 VDD!  PFET  L=200E-9 W=4.1E-6 AD=+2.05000000E-12 
+AS=+2.05000000E-12 PD=+9.20000000E-06 PS=+9.20000000E-06 NRD=+1.21951220E-01 
+NRS=+1.21951220E-01 M=1.0 
M31 RDECO_7 RIB_0 NET062 VDD!  PFET  L=200E-9 W=4.1E-6 AD=+2.05000000E-12 
+AS=+2.05000000E-12 PD=+9.20000000E-06 PS=+9.20000000E-06 NRD=+1.21951220E-01 
+NRS=+1.21951220E-01 M=1.0 
M8 RDECO_0 RI_0 NET056 VDD!  PFET  L=200E-9 W=4.1E-6 AD=+2.05000000E-12 
+AS=+2.05000000E-12 PD=+9.20000000E-06 PS=+9.20000000E-06 NRD=+1.21951220E-01 
+NRS=+1.21951220E-01 M=1.0 
M27 RDECO_6 RI_0 NET062 VDD!  PFET  L=200E-9 W=4.1E-6 AD=+2.05000000E-12 
+AS=+2.05000000E-12 PD=+9.20000000E-06 PS=+9.20000000E-06 NRD=+1.21951220E-01 
+NRS=+1.21951220E-01 M=1.0 
M32 NET056 RI_1 NET0175 VDD!  PFET  L=200E-9 W=8.2E-6 AD=+4.10000000E-12 
+AS=+4.10000000E-12 PD=+1.74000000E-05 PS=+1.74000000E-05 NRD=+6.09756098E-02 
+NRS=+6.09756098E-02 M=1.0 
M33 NET050 RI_1 NET0174 VDD!  PFET  L=200E-9 W=8.2E-6 AD=+4.10000000E-12 
+AS=+4.10000000E-12 PD=+1.74000000E-05 PS=+1.74000000E-05 NRD=+6.09756098E-02 
+NRS=+6.09756098E-02 M=1.0 
M34 NET068 RIB_1 NET0175 VDD!  PFET  L=200E-9 W=8.2E-6 AD=+4.10000000E-12 
+AS=+4.10000000E-12 PD=+1.74000000E-05 PS=+1.74000000E-05 NRD=+6.09756098E-02 
+NRS=+6.09756098E-02 M=1.0 
M35 NET062 RIB_1 NET0174 VDD!  PFET  L=200E-9 W=8.2E-6 AD=+4.10000000E-12 
+AS=+4.10000000E-12 PD=+1.74000000E-05 PS=+1.74000000E-05 NRD=+6.09756098E-02 
+NRS=+6.09756098E-02 M=1.0 
M26 RDECO_4 RI_0 NET050 VDD!  PFET  L=200E-9 W=4.1E-6 AD=+2.05000000E-12 
+AS=+2.05000000E-12 PD=+9.20000000E-06 PS=+9.20000000E-06 NRD=+1.21951220E-01 
+NRS=+1.21951220E-01 M=1.0 
M25 RDECO_2 RI_0 NET068 VDD!  PFET  L=200E-9 W=4.1E-6 AD=+2.05000000E-12 
+AS=+2.05000000E-12 PD=+9.20000000E-06 PS=+9.20000000E-06 NRD=+1.21951220E-01 
+NRS=+1.21951220E-01 M=1.0 
M24 RDECO_0 RI_1 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M23 RDECO_7 RIB_2 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M22 RDECO_6 RIB_2 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M21 RDECO_5 RIB_2 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M20 RDECO_4 RIB_2 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M19 RDECO_3 RI_2 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M18 RDECO_2 RI_2 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M17 RDECO_1 RI_2 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M16 RDECO_0 RI_2 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M15 RDECO_7 RIB_1 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M14 RDECO_6 RIB_1 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M13 RDECO_3 RIB_1 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M12 RDECO_2 RIB_1 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M11 RDECO_5 RI_1 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M10 RDECO_4 RI_1 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M9 RDECO_1 RI_1 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M7 RDECO_7 RIB_0 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M6 RDECO_5 RIB_0 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M5 RDECO_3 RIB_0 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M4 RDECO_1 RIB_0 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M3 RDECO_6 RI_0 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M2 RDECO_4 RI_0 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M1 RDECO_2 RI_0 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M0 RDECO_0 RI_0 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS RDEC3TO8A_G7 
* FILE NAME: SRAM2_SAMP_CELL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SAMP_CELL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:43 2007.
   
* TERMINAL MAPPING: BIT = BIT
*                   OUT = OUT
*                   BIT_BAR = BIT_BAR
*                   OUT_BAR = OUT_BAR
*                   SENSE_DISABLE = SENSE_DISABLE
.SUBCKT SAMP_CELL_G12 BIT OUT BIT_BAR OUT_BAR SENSE_DISABLE 
M4 OUT OUT_BAR VDD! VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M3 OUT_BAR OUT VDD! VDD!  PFET  L=200E-9 W=400E-9 AD=+2.00000000E-13 
+AS=+2.00000000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 NRD=+1.25000000E+00 
+NRS=+1.25000000E+00 M=1.0 
M2 OUT_BAR SENSE_DISABLE BIT_BAR VDD!  PFET  L=200E-9 W=3.6E-6 
+AD=+1.80000000E-12 AS=+1.80000000E-12 PD=+8.20000000E-06 PS=+8.20000000E-06 
+NRD=+1.38888889E-01 NRS=+1.38888889E-01 M=1.0 
M1 OUT SENSE_DISABLE BIT VDD!  PFET  L=200E-9 W=3.6E-6 AD=+1.80000000E-12 
+AS=+1.80000000E-12 PD=+8.20000000E-06 PS=+8.20000000E-06 NRD=+1.38888889E-01 
+NRS=+1.38888889E-01 M=1.0 
M6 OUT OUT_BAR NET20 0  NFET  L=200E-9 W=3.6E-6 AD=+1.80000000E-12 
+AS=+1.80000000E-12 PD=+8.20000000E-06 PS=+8.20000000E-06 NRD=+1.38888889E-01 
+NRS=+1.38888889E-01 M=1.0 
M5 OUT_BAR OUT NET20 0  NFET  L=200E-9 W=3.6E-6 AD=+1.80000000E-12 
+AS=+1.80000000E-12 PD=+8.20000000E-06 PS=+8.20000000E-06 NRD=+1.38888889E-01 
+NRS=+1.38888889E-01 M=1.0 
M0 NET20 SENSE_DISABLE 0 0  NFET  L=200E-9 W=3.6E-6 AD=+1.80000000E-12 
+AS=+1.80000000E-12 PD=+8.20000000E-06 PS=+8.20000000E-06 NRD=+1.38888889E-01 
+NRS=+1.38888889E-01 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SAMP_CELL_G12 
* FILE NAME: SRAM2_SRAM_CELL64X32_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SRAM_CELL64X32.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:40 2007.
   
* TERMINAL MAPPING: BIT<0> = BIT_0
*                   BIT<1> = BIT_1
*                   BIT<2> = BIT_2
*                   BIT<3> = BIT_3
*                   BIT<4> = BIT_4
*                   BIT<5> = BIT_5
*                   BIT<6> = BIT_6
*                   BIT<7> = BIT_7
*                   BIT<8> = BIT_8
*                   BIT<9> = BIT_9
*                   BIT<10> = BIT_10
*                   BIT<11> = BIT_11
*                   BIT<12> = BIT_12
*                   BIT<13> = BIT_13
*                   BIT<14> = BIT_14
*                   BIT<15> = BIT_15
*                   BIT<16> = BIT_16
*                   BIT<17> = BIT_17
*                   BIT<18> = BIT_18
*                   BIT<19> = BIT_19
*                   BIT<20> = BIT_20
*                   BIT<21> = BIT_21
*                   BIT<22> = BIT_22
*                   BIT<23> = BIT_23
*                   BIT<24> = BIT_24
*                   BIT<25> = BIT_25
*                   BIT<26> = BIT_26
*                   BIT<27> = BIT_27
*                   BIT<28> = BIT_28
*                   BIT<29> = BIT_29
*                   BIT<30> = BIT_30
*                   BIT<31> = BIT_31
*                   BIT_B<0> = BIT_B_0
*                   BIT_B<1> = BIT_B_1
*                   BIT_B<2> = BIT_B_2
*                   BIT_B<3> = BIT_B_3
*                   BIT_B<4> = BIT_B_4
*                   BIT_B<5> = BIT_B_5
*                   BIT_B<6> = BIT_B_6
*                   BIT_B<7> = BIT_B_7
*                   BIT_B<8> = BIT_B_8
*                   BIT_B<9> = BIT_B_9
*                   BIT_B<10> = BIT_B_10
*                   BIT_B<11> = BIT_B_11
*                   BIT_B<12> = BIT_B_12
*                   BIT_B<13> = BIT_B_13
*                   BIT_B<14> = BIT_B_14
*                   BIT_B<15> = BIT_B_15
*                   BIT_B<16> = BIT_B_16
*                   BIT_B<17> = BIT_B_17
*                   BIT_B<18> = BIT_B_18
*                   BIT_B<19> = BIT_B_19
*                   BIT_B<20> = BIT_B_20
*                   BIT_B<21> = BIT_B_21
*                   BIT_B<22> = BIT_B_22
*                   BIT_B<23> = BIT_B_23
*                   BIT_B<24> = BIT_B_24
*                   BIT_B<25> = BIT_B_25
*                   BIT_B<26> = BIT_B_26
*                   BIT_B<27> = BIT_B_27
*                   BIT_B<28> = BIT_B_28
*                   BIT_B<29> = BIT_B_29
*                   BIT_B<30> = BIT_B_30
*                   BIT_B<31> = BIT_B_31
*                   WL<0> = WL_0
*                   WL<1> = WL_1
*                   WL<2> = WL_2
*                   WL<3> = WL_3
*                   WL<4> = WL_4
*                   WL<5> = WL_5
*                   WL<6> = WL_6
*                   WL<7> = WL_7
*                   WL<8> = WL_8
*                   WL<9> = WL_9
*                   WL<10> = WL_10
*                   WL<11> = WL_11
*                   WL<12> = WL_12
*                   WL<13> = WL_13
*                   WL<14> = WL_14
*                   WL<15> = WL_15
*                   WL<16> = WL_16
*                   WL<17> = WL_17
*                   WL<18> = WL_18
*                   WL<19> = WL_19
*                   WL<20> = WL_20
*                   WL<21> = WL_21
*                   WL<22> = WL_22
*                   WL<23> = WL_23
*                   WL<24> = WL_24
*                   WL<25> = WL_25
*                   WL<26> = WL_26
*                   WL<27> = WL_27
*                   WL<28> = WL_28
*                   WL<29> = WL_29
*                   WL<30> = WL_30
*                   WL<31> = WL_31
*                   WL<32> = WL_32
*                   WL<33> = WL_33
*                   WL<34> = WL_34
*                   WL<35> = WL_35
*                   WL<36> = WL_36
*                   WL<37> = WL_37
*                   WL<38> = WL_38
*                   WL<39> = WL_39
*                   WL<40> = WL_40
*                   WL<41> = WL_41
*                   WL<42> = WL_42
*                   WL<43> = WL_43
*                   WL<44> = WL_44
*                   WL<45> = WL_45
*                   WL<46> = WL_46
*                   WL<47> = WL_47
*                   WL<48> = WL_48
*                   WL<49> = WL_49
*                   WL<50> = WL_50
*                   WL<51> = WL_51
*                   WL<52> = WL_52
*                   WL<53> = WL_53
*                   WL<54> = WL_54
*                   WL<55> = WL_55
*                   WL<56> = WL_56
*                   WL<57> = WL_57
*                   WL<58> = WL_58
*                   WL<59> = WL_59
*                   WL<60> = WL_60
*                   WL<61> = WL_61
*                   WL<62> = WL_62
*                   WL<63> = WL_63
.SUBCKT SUB2 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 BIT_8 BIT_9 
+BIT_10 BIT_11 BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 BIT_19 BIT_20 
+BIT_21 BIT_22 BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 BIT_30 BIT_31 
+BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 BIT_B_4 BIT_B_5 BIT_B_6 BIT_B_7 BIT_B_8 
+BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 BIT_B_13 BIT_B_14 BIT_B_15 BIT_B_16 
+BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 BIT_B_21 BIT_B_22 BIT_B_23 BIT_B_24 
+BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 BIT_B_29 BIT_B_30 BIT_B_31 WL_0 WL_1 WL_2 
+WL_3 WL_4 WL_5 WL_6 WL_7 WL_8 WL_9 WL_10 WL_11 WL_12 WL_13 WL_14 WL_15 WL_16 
+WL_17 WL_18 WL_19 WL_20 WL_21 WL_22 WL_23 WL_24 WL_25 WL_26 WL_27 WL_28 WL_29 
+WL_30 WL_31 WL_32 WL_33 WL_34 WL_35 WL_36 WL_37 WL_38 WL_39 WL_40 WL_41 WL_42 
+WL_43 WL_44 WL_45 WL_46 WL_47 WL_48 WL_49 WL_50 WL_51 WL_52 WL_53 WL_54 WL_55 
+WL_56 WL_57 WL_58 WL_59 WL_60 WL_61 WL_62 WL_63 
XI65 BIT_0 BIT_1 BIT_2 BIT_3 BIT_4 BIT_5 BIT_6 BIT_7 BIT_8 BIT_9 BIT_10 BIT_11 
+BIT_12 BIT_13 BIT_14 BIT_15 BIT_16 BIT_17 BIT_18 BIT_19 BIT_20 BIT_21 BIT_22 
+BIT_23 BIT_24 BIT_25 BIT_26 BIT_27 BIT_28 BIT_29 BIT_30 BIT_31 NET201_0 
+NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 NET201_8 
+NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 NET201_16 
+NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 NET201_23 
+NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 NET201_30 
+NET201_31 TL_PI_MODEL32_1 
XI66 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 NET203_6 NET203_7 
+NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 NET203_14 NET203_15 
+NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 NET203_21 NET203_22 
+NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 NET203_28 NET203_29 
+NET203_30 NET203_31 BIT_B_0 BIT_B_1 BIT_B_2 BIT_B_3 BIT_B_4 BIT_B_5 BIT_B_6 
+BIT_B_7 BIT_B_8 BIT_B_9 BIT_B_10 BIT_B_11 BIT_B_12 BIT_B_13 BIT_B_14 BIT_B_15 
+BIT_B_16 BIT_B_17 BIT_B_18 BIT_B_19 BIT_B_20 BIT_B_21 BIT_B_22 BIT_B_23 
+BIT_B_24 BIT_B_25 BIT_B_26 BIT_B_27 BIT_B_28 BIT_B_29 BIT_B_30 BIT_B_31 
+TL_PI_MODEL32_1 
XI63 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_63 SRAM_CELL32_G3 
XI62 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_62 SRAM_CELL32_G3 
XI61 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_61 SRAM_CELL32_G3 
XI60 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_60 SRAM_CELL32_G3 
XI59 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_59 SRAM_CELL32_G3 
XI58 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_58 SRAM_CELL32_G3 
XI57 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_57 SRAM_CELL32_G3 
XI56 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_56 SRAM_CELL32_G3 
XI55 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_55 SRAM_CELL32_G3 
XI54 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_54 SRAM_CELL32_G3 
XI53 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_53 SRAM_CELL32_G3 
XI52 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_52 SRAM_CELL32_G3 
XI51 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_51 SRAM_CELL32_G3 
XI50 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_50 SRAM_CELL32_G3 
XI49 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_49 SRAM_CELL32_G3 
XI48 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_48 SRAM_CELL32_G3 
XI47 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_47 SRAM_CELL32_G3 
XI46 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_46 SRAM_CELL32_G3 
XI45 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_45 SRAM_CELL32_G3 
XI44 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_44 SRAM_CELL32_G3 
XI43 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_43 SRAM_CELL32_G3 
XI42 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_42 SRAM_CELL32_G3 
XI41 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_41 SRAM_CELL32_G3 
XI40 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_40 SRAM_CELL32_G3 
XI39 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_39 SRAM_CELL32_G3 
XI38 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_38 SRAM_CELL32_G3 
XI37 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_37 SRAM_CELL32_G3 
XI36 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_36 SRAM_CELL32_G3 
XI35 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_35 SRAM_CELL32_G3 
XI34 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_34 SRAM_CELL32_G3 
XI33 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_33 SRAM_CELL32_G3 
XI32 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_32 SRAM_CELL32_G3 
XI31 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_31 SRAM_CELL32_G3 
XI30 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_30 SRAM_CELL32_G3 
XI29 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_29 SRAM_CELL32_G3 
XI28 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_28 SRAM_CELL32_G3 
XI27 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_27 SRAM_CELL32_G3 
XI26 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_26 SRAM_CELL32_G3 
XI25 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_25 SRAM_CELL32_G3 
XI24 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_24 SRAM_CELL32_G3 
XI23 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_23 SRAM_CELL32_G3 
XI22 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_22 SRAM_CELL32_G3 
XI21 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_21 SRAM_CELL32_G3 
XI20 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_20 SRAM_CELL32_G3 
XI19 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_19 SRAM_CELL32_G3 
XI18 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_18 SRAM_CELL32_G3 
XI17 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_17 SRAM_CELL32_G3 
XI16 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_16 SRAM_CELL32_G3 
XI15 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_15 SRAM_CELL32_G3 
XI14 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_14 SRAM_CELL32_G3 
XI13 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_13 SRAM_CELL32_G3 
XI12 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_12 SRAM_CELL32_G3 
XI11 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_11 SRAM_CELL32_G3 
XI10 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_10 SRAM_CELL32_G3 
XI9 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_9 SRAM_CELL32_G3 
XI8 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_8 SRAM_CELL32_G3 
XI7 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_7 SRAM_CELL32_G3 
XI6 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_6 SRAM_CELL32_G3 
XI5 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_5 SRAM_CELL32_G3 
XI4 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_4 SRAM_CELL32_G3 
XI3 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_3 SRAM_CELL32_G3 
XI2 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_2 SRAM_CELL32_G3 
XI1 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_1 SRAM_CELL32_G3 
XI0 NET201_0 NET201_1 NET201_2 NET201_3 NET201_4 NET201_5 NET201_6 NET201_7 
+NET201_8 NET201_9 NET201_10 NET201_11 NET201_12 NET201_13 NET201_14 NET201_15 
+NET201_16 NET201_17 NET201_18 NET201_19 NET201_20 NET201_21 NET201_22 
+NET201_23 NET201_24 NET201_25 NET201_26 NET201_27 NET201_28 NET201_29 
+NET201_30 NET201_31 NET203_0 NET203_1 NET203_2 NET203_3 NET203_4 NET203_5 
+NET203_6 NET203_7 NET203_8 NET203_9 NET203_10 NET203_11 NET203_12 NET203_13 
+NET203_14 NET203_15 NET203_16 NET203_17 NET203_18 NET203_19 NET203_20 
+NET203_21 NET203_22 NET203_23 NET203_24 NET203_25 NET203_26 NET203_27 
+NET203_28 NET203_29 NET203_30 NET203_31 WL_0 SRAM_CELL32_G3 
   
   
* FILE NAME: SRAM2_TL_PI_MODEL32_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL32.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:32 2007.
   
* TERMINAL MAPPING: IN<0> = IN_0
*                   IN<1> = IN_1
*                   IN<2> = IN_2
*                   IN<3> = IN_3
*                   IN<4> = IN_4
*                   IN<5> = IN_5
*                   IN<6> = IN_6
*                   IN<7> = IN_7
*                   IN<8> = IN_8
*                   IN<9> = IN_9
*                   IN<10> = IN_10
*                   IN<11> = IN_11
*                   IN<12> = IN_12
*                   IN<13> = IN_13
*                   IN<14> = IN_14
*                   IN<15> = IN_15
*                   IN<16> = IN_16
*                   IN<17> = IN_17
*                   IN<18> = IN_18
*                   IN<19> = IN_19
*                   IN<20> = IN_20
*                   IN<21> = IN_21
*                   IN<22> = IN_22
*                   IN<23> = IN_23
*                   IN<24> = IN_24
*                   IN<25> = IN_25
*                   IN<26> = IN_26
*                   IN<27> = IN_27
*                   IN<28> = IN_28
*                   IN<29> = IN_29
*                   IN<30> = IN_30
*                   IN<31> = IN_31
*                   OUT<0> = OUT_0
*                   OUT<1> = OUT_1
*                   OUT<2> = OUT_2
*                   OUT<3> = OUT_3
*                   OUT<4> = OUT_4
*                   OUT<5> = OUT_5
*                   OUT<6> = OUT_6
*                   OUT<7> = OUT_7
*                   OUT<8> = OUT_8
*                   OUT<9> = OUT_9
*                   OUT<10> = OUT_10
*                   OUT<11> = OUT_11
*                   OUT<12> = OUT_12
*                   OUT<13> = OUT_13
*                   OUT<14> = OUT_14
*                   OUT<15> = OUT_15
*                   OUT<16> = OUT_16
*                   OUT<17> = OUT_17
*                   OUT<18> = OUT_18
*                   OUT<19> = OUT_19
*                   OUT<20> = OUT_20
*                   OUT<21> = OUT_21
*                   OUT<22> = OUT_22
*                   OUT<23> = OUT_23
*                   OUT<24> = OUT_24
*                   OUT<25> = OUT_25
*                   OUT<26> = OUT_26
*                   OUT<27> = OUT_27
*                   OUT<28> = OUT_28
*                   OUT<29> = OUT_29
*                   OUT<30> = OUT_30
*                   OUT<31> = OUT_31
.SUBCKT TL_PI_MODEL32_1 IN_0 IN_1 IN_2 IN_3 IN_4 IN_5 IN_6 IN_7 IN_8 IN_9 
+IN_10 IN_11 IN_12 IN_13 IN_14 IN_15 IN_16 IN_17 IN_18 IN_19 IN_20 IN_21 IN_22 
+IN_23 IN_24 IN_25 IN_26 IN_27 IN_28 IN_29 IN_30 IN_31 OUT_0 OUT_1 OUT_2 OUT_3 
+OUT_4 OUT_5 OUT_6 OUT_7 OUT_8 OUT_9 OUT_10 OUT_11 OUT_12 OUT_13 OUT_14 OUT_15 
+OUT_16 OUT_17 OUT_18 OUT_19 OUT_20 OUT_21 OUT_22 OUT_23 OUT_24 OUT_25 OUT_26 
+OUT_27 OUT_28 OUT_29 OUT_30 OUT_31 
XI31 IN_31 OUT_31 TL_PI_MODEL_1 
XI30 IN_30 OUT_30 TL_PI_MODEL_1 
XI29 IN_29 OUT_29 TL_PI_MODEL_1 
XI28 IN_28 OUT_28 TL_PI_MODEL_1 
XI27 IN_27 OUT_27 TL_PI_MODEL_1 
XI26 IN_26 OUT_26 TL_PI_MODEL_1 
XI25 IN_25 OUT_25 TL_PI_MODEL_1 
XI24 IN_24 OUT_24 TL_PI_MODEL_1 
XI23 IN_23 OUT_23 TL_PI_MODEL_1 
XI22 IN_22 OUT_22 TL_PI_MODEL_1 
XI21 IN_21 OUT_21 TL_PI_MODEL_1 
XI20 IN_20 OUT_20 TL_PI_MODEL_1 
XI19 IN_19 OUT_19 TL_PI_MODEL_1 
XI18 IN_18 OUT_18 TL_PI_MODEL_1 
XI17 IN_17 OUT_17 TL_PI_MODEL_1 
XI16 IN_16 OUT_16 TL_PI_MODEL_1 
XI15 IN_15 OUT_15 TL_PI_MODEL_1 
XI14 IN_14 OUT_14 TL_PI_MODEL_1 
XI13 IN_13 OUT_13 TL_PI_MODEL_1 
XI12 IN_12 OUT_12 TL_PI_MODEL_1 
XI11 IN_11 OUT_11 TL_PI_MODEL_1 
XI10 IN_10 OUT_10 TL_PI_MODEL_1 
XI9 IN_9 OUT_9 TL_PI_MODEL_1 
XI8 IN_8 OUT_8 TL_PI_MODEL_1 
XI7 IN_7 OUT_7 TL_PI_MODEL_1 
XI6 IN_6 OUT_6 TL_PI_MODEL_1 
XI5 IN_5 OUT_5 TL_PI_MODEL_1 
XI4 IN_4 OUT_4 TL_PI_MODEL_1 
XI3 IN_3 OUT_3 TL_PI_MODEL_1 
XI2 IN_2 OUT_2 TL_PI_MODEL_1 
XI1 IN_1 OUT_1 TL_PI_MODEL_1 
XI0 IN_0 OUT_0 TL_PI_MODEL_1 
   
   
* FILE NAME: SRAM2_TL_PI_MODEL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TL_PI_MODEL.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:31 2007.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT TL_PI_MODEL_1 IN OUT 
C0 IN 0  ((33.8E-15)) M=1.0 
C1 OUT 0  ((33.8E-15)) M=1.0 
R0 IN OUT  ((179.2)) M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TL_PI_MODEL32_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SUB2 
* FILE NAME: SRAM_RDEC4TO16A_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: RDEC4TO16A.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:38 2007.
   
* TERMINAL MAPPING: RDECO<0> = RDECO_0
*                   RDECO<1> = RDECO_1
*                   RDECO<2> = RDECO_2
*                   RDECO<3> = RDECO_3
*                   RDECO<4> = RDECO_4
*                   RDECO<5> = RDECO_5
*                   RDECO<6> = RDECO_6
*                   RDECO<7> = RDECO_7
*                   RDECO<8> = RDECO_8
*                   RDECO<9> = RDECO_9
*                   RDECO<10> = RDECO_10
*                   RDECO<11> = RDECO_11
*                   RDECO<12> = RDECO_12
*                   RDECO<13> = RDECO_13
*                   RDECO<14> = RDECO_14
*                   RDECO<15> = RDECO_15
*                   RI<0> = RI_0
*                   RI<1> = RI_1
*                   RI<2> = RI_2
*                   RI<3> = RI_3
*                   RIB<0> = RIB_0
*                   RIB<1> = RIB_1
*                   RIB<2> = RIB_2
*                   RIB<3> = RIB_3
*                   TOP = TOP
.SUBCKT RDEC4TO16A_G8 RDECO_0 RDECO_1 RDECO_2 RDECO_3 RDECO_4 RDECO_5 RDECO_6 
+RDECO_7 RDECO_8 RDECO_9 RDECO_10 RDECO_11 RDECO_12 RDECO_13 RDECO_14 RDECO_15 
+RI_0 RI_1 RI_2 RI_3 RIB_0 RIB_1 RIB_2 RIB_3 TOP 
XI8 RDECO_0 RDECO_1 RDECO_2 RDECO_3 RDECO_4 RDECO_5 RDECO_6 RDECO_7 RI_0 RI_1 
+RI_2 RIB_0 RIB_1 RIB_2 NET75 RDEC3TO8A_G7 
XI9 RDECO_8 RDECO_9 RDECO_10 RDECO_11 RDECO_12 RDECO_13 RDECO_14 RDECO_15 RI_0 
+RI_1 RI_2 RIB_0 RIB_1 RIB_2 NET90 RDEC3TO8A_G7 
M12 RDECO_14 RIB_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M13 RDECO_13 RIB_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M11 RDECO_15 RIB_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M14 RDECO_12 RIB_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M15 RDECO_11 RIB_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M16 RDECO_10 RIB_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M17 RDECO_9 RIB_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M18 RDECO_8 RIB_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M2 RDECO_7 RI_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M3 RDECO_6 RI_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M4 RDECO_5 RI_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M5 RDECO_4 RI_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M6 RDECO_3 RI_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M7 RDECO_2 RI_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M8 RDECO_1 RI_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M9 RDECO_0 RI_3 0 0  NFET  L=200E-9 W=1.4E-6 AD=+7.00000000E-13 
+AS=+7.00000000E-13 PD=+3.80000000E-06 PS=+3.80000000E-06 NRD=+3.57142857E-01 
+NRS=+3.57142857E-01 M=1.0 
M1 NET90 RIB_3 TOP VDD!  PFET  L=200E-9 W=36.8E-6 AD=+1.84000000E-11 
+AS=+1.84000000E-11 PD=+7.46000000E-05 PS=+7.46000000E-05 NRD=+1.35869565E-02 
+NRS=+1.35869565E-02 M=1.0 
M0 NET75 RI_3 TOP VDD!  PFET  L=200E-9 W=36.8E-6 AD=+1.84000000E-11 
+AS=+1.84000000E-11 PD=+7.46000000E-05 PS=+7.46000000E-05 NRD=+1.35869565E-02 
+NRS=+1.35869565E-02 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS RDEC4TO16A_G8 
* FILE NAME: OSU_STDCELLS_CLKBUF3_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: CLKBUF3.
* GENERATED FOR: HSPICES.
* GENERATED ON OCT 25 01:12:33 2007.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT CLKBUF3_G16 A Y 
M8 NET145 NET142 VDD! VDD!  TSMC20P  L=200E-9 W=8E-6 AD=4E-12 AS=4E-12 
+PD=17E-6 PS=17E-6 M=1 
M9 NET142 NET139 VDD! VDD!  TSMC20P  L=200E-9 W=8E-6 AD=4E-12 AS=4E-12 
+PD=17E-6 PS=17E-6 M=1 
M10 NET139 NET136 VDD! VDD!  TSMC20P  L=200E-9 W=8E-6 AD=4E-12 AS=4E-12 
+PD=17E-6 PS=17E-6 M=1 
M11 NET136 A VDD! VDD!  TSMC20P  L=200E-9 W=8E-6 AD=4E-12 AS=4E-12 PD=17E-6 
+PS=17E-6 M=1 
M0 NET157 NET145 VDD! VDD!  TSMC20P  L=200E-9 W=8E-6 AD=4E-12 AS=4E-12 
+PD=17E-6 PS=17E-6 M=1 
M3 NET154 NET157 VDD! VDD!  TSMC20P  L=200E-9 W=8E-6 AD=4E-12 AS=4E-12 
+PD=17E-6 PS=17E-6 M=1 
M5 NET151 NET154 VDD! VDD!  TSMC20P  L=200E-9 W=8E-6 AD=4E-12 AS=4E-12 
+PD=17E-6 PS=17E-6 M=1 
M6 Y NET151 VDD! VDD!  TSMC20P  L=200E-9 W=8E-6 AD=4E-12 AS=4E-12 PD=17E-6 
+PS=17E-6 M=1 
M12 NET145 NET142 0 0  TSMC20N  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M13 NET142 NET139 0 0  TSMC20N  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M14 NET139 NET136 0 0  TSMC20N  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M15 NET136 A 0 0  TSMC20N  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 PS=9E-6 
+M=1 
M1 NET157 NET145 0 0  TSMC20N  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M2 NET154 NET157 0 0  TSMC20N  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M4 NET151 NET154 0 0  TSMC20N  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M7 Y NET151 0 0  TSMC20N  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 PS=9E-6 
+M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS CLKBUF3_G16 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc20P" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc20N" NMOS 
   
   
* INCLUDE FILES
   
   
   
   
   
   
* END OF NETLIST
.TEMP    75.0000    
.OP
.save
.OPTION  INGOLD=2 ARTIST=2 PSF=2
+        PROBE=0
.END
